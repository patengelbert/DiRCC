// dircc_avalon_st_packet_sender_tb.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_avalon_st_packet_sender_tb (
	);

	import dircc_types_pkg::*;

	wire         dircc_avalon_st_packet_sender_inst_output_valid;                 
	wire  [31:0] dircc_avalon_st_packet_sender_inst_output_data;                  
	wire         dircc_avalon_st_packet_sender_inst_output_ready;                 
	wire         dircc_avalon_st_packet_sender_inst_output_startofpacket;         
	wire         dircc_avalon_st_packet_sender_inst_output_endofpacket;           
	wire   [1:0] dircc_avalon_st_packet_sender_inst_output_empty;
	wire         dircc_avalon_st_packet_sender_inst_clk_bfm_clk_clk;
	wire         dircc_avalon_st_packet_sender_inst_reset_bfm_reset_reset;
	wire         dircc_avalon_st_packet_sender_inst_sending;
	packet_t	 dircc_avalon_st_packet_sender_inst_packet_data;
	logic 		 dircc_avalon_st_packet_sender_inst_write_packet;

	dircc_avalon_st_packet_sender dircc_avalon_st_packet_sender_inst (
		.clk	                    (dircc_avalon_st_packet_sender_inst_clk_bfm_clk_clk),                   //          clk.clk
		.data           			(dircc_avalon_st_packet_sender_inst_output_data),                  		//  	 output.data
		.valid          			(dircc_avalon_st_packet_sender_inst_output_valid),                 		//             .valid
		.ready          			(dircc_avalon_st_packet_sender_inst_output_ready),                 		//             .ready
		.startofpacket  			(dircc_avalon_st_packet_sender_inst_output_startofpacket),         		//             .startofpacket
		.endofpacket    			(dircc_avalon_st_packet_sender_inst_output_endofpacket),           		//             .endofpacket
		.empty          			(dircc_avalon_st_packet_sender_inst_output_empty),                 		//             .empty
		.reset_n              		(dircc_avalon_st_packet_sender_inst_reset_bfm_reset_reset),             //        reset.reset_n
		.sending					(dircc_avalon_st_packet_sender_inst_sending),							//		sending.sending
		.packet_data				(dircc_avalon_st_packet_sender_inst_packet_data),						//		 packet.data
		.write_packet				(dircc_avalon_st_packet_sender_inst_write_packet)						//		   	   .write_packet
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dircc_avalon_st_packet_sender_inst_clk_bfm (
		.clk (dircc_avalon_st_packet_sender_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dircc_avalon_st_packet_sender_inst_output_bfm (
		.clk                (dircc_avalon_st_packet_sender_inst_clk_bfm_clk_clk),           //       clk.clk
		.reset              (~dircc_avalon_st_packet_sender_inst_reset_bfm_reset_reset),    // clk_reset.reset
		.sink_data          (dircc_avalon_st_packet_sender_inst_output_data),          		//      sink.data
		.sink_valid         (dircc_avalon_st_packet_sender_inst_output_valid),         		//          .valid
		.sink_ready         (dircc_avalon_st_packet_sender_inst_output_ready),         		//          .ready
		.sink_startofpacket (dircc_avalon_st_packet_sender_inst_output_startofpacket), 		//          .startofpacket
		.sink_endofpacket   (dircc_avalon_st_packet_sender_inst_output_endofpacket),   		//          .endofpacket
		.sink_empty         (dircc_avalon_st_packet_sender_inst_output_empty),         		//          .empty
		.sink_channel       (1'b0),                                         				// (terminated)
		.sink_error         (1'b0)                                          				// (terminated)
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dircc_avalon_st_packet_sender_inst_reset_bfm (
		.reset (dircc_avalon_st_packet_sender_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dircc_avalon_st_packet_sender_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
