// dircc_routing_tb.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_routing_tb (
	);

	wire         dircc_routing_inst_output_east_valid;                 // dircc_routing_inst:output_east_valid -> dircc_routing_inst_output_east_bfm:sink_valid
	wire  [31:0] dircc_routing_inst_output_east_data;                  // dircc_routing_inst:output_east_data -> dircc_routing_inst_output_east_bfm:sink_data
	wire         dircc_routing_inst_output_east_ready;                 // dircc_routing_inst_output_east_bfm:sink_ready -> dircc_routing_inst:output_east_ready
	wire         dircc_routing_inst_output_east_startofpacket;         // dircc_routing_inst:output_east_startofpacket -> dircc_routing_inst_output_east_bfm:sink_startofpacket
	wire         dircc_routing_inst_output_east_endofpacket;           // dircc_routing_inst:output_east_endofpacket -> dircc_routing_inst_output_east_bfm:sink_endofpacket
	wire   [1:0] dircc_routing_inst_output_east_empty;                 // dircc_routing_inst:output_east_empty -> dircc_routing_inst_output_east_bfm:sink_empty
	wire         dircc_routing_inst_output_here_valid;                 // dircc_routing_inst:output_here_valid -> dircc_routing_inst_output_here_bfm:sink_valid
	wire  [31:0] dircc_routing_inst_output_here_data;                  // dircc_routing_inst:output_here_data -> dircc_routing_inst_output_here_bfm:sink_data
	wire         dircc_routing_inst_output_here_ready;                 // dircc_routing_inst_output_here_bfm:sink_ready -> dircc_routing_inst:output_here_ready
	wire         dircc_routing_inst_output_here_startofpacket;         // dircc_routing_inst:output_here_startofpacket -> dircc_routing_inst_output_here_bfm:sink_startofpacket
	wire         dircc_routing_inst_output_here_endofpacket;           // dircc_routing_inst:output_here_endofpacket -> dircc_routing_inst_output_here_bfm:sink_endofpacket
	wire   [1:0] dircc_routing_inst_output_here_empty;                 // dircc_routing_inst:output_here_empty -> dircc_routing_inst_output_here_bfm:sink_empty
	wire         dircc_routing_inst_output_north_valid;                // dircc_routing_inst:output_north_valid -> dircc_routing_inst_output_north_bfm:sink_valid
	wire  [31:0] dircc_routing_inst_output_north_data;                 // dircc_routing_inst:output_north_data -> dircc_routing_inst_output_north_bfm:sink_data
	wire         dircc_routing_inst_output_north_ready;                // dircc_routing_inst_output_north_bfm:sink_ready -> dircc_routing_inst:output_north_ready
	wire         dircc_routing_inst_output_north_startofpacket;        // dircc_routing_inst:output_north_startofpacket -> dircc_routing_inst_output_north_bfm:sink_startofpacket
	wire         dircc_routing_inst_output_north_endofpacket;          // dircc_routing_inst:output_north_endofpacket -> dircc_routing_inst_output_north_bfm:sink_endofpacket
	wire   [1:0] dircc_routing_inst_output_north_empty;                // dircc_routing_inst:output_north_empty -> dircc_routing_inst_output_north_bfm:sink_empty
	wire         dircc_routing_inst_output_south_valid;                // dircc_routing_inst:output_south_valid -> dircc_routing_inst_output_south_bfm:sink_valid
	wire  [31:0] dircc_routing_inst_output_south_data;                 // dircc_routing_inst:output_south_data -> dircc_routing_inst_output_south_bfm:sink_data
	wire         dircc_routing_inst_output_south_ready;                // dircc_routing_inst_output_south_bfm:sink_ready -> dircc_routing_inst:output_south_ready
	wire         dircc_routing_inst_output_south_startofpacket;        // dircc_routing_inst:output_south_startofpacket -> dircc_routing_inst_output_south_bfm:sink_startofpacket
	wire         dircc_routing_inst_output_south_endofpacket;          // dircc_routing_inst:output_south_endofpacket -> dircc_routing_inst_output_south_bfm:sink_endofpacket
	wire   [1:0] dircc_routing_inst_output_south_empty;                // dircc_routing_inst:output_south_empty -> dircc_routing_inst_output_south_bfm:sink_empty
	wire         dircc_routing_inst_output_west_valid;                 // dircc_routing_inst:output_west_valid -> dircc_routing_inst_output_west_bfm:sink_valid
	wire  [31:0] dircc_routing_inst_output_west_data;                  // dircc_routing_inst:output_west_data -> dircc_routing_inst_output_west_bfm:sink_data
	wire         dircc_routing_inst_output_west_ready;                 // dircc_routing_inst_output_west_bfm:sink_ready -> dircc_routing_inst:output_west_ready
	wire         dircc_routing_inst_output_west_startofpacket;         // dircc_routing_inst:output_west_startofpacket -> dircc_routing_inst_output_west_bfm:sink_startofpacket
	wire         dircc_routing_inst_output_west_endofpacket;           // dircc_routing_inst:output_west_endofpacket -> dircc_routing_inst_output_west_bfm:sink_endofpacket
	wire   [1:0] dircc_routing_inst_output_west_empty;                 // dircc_routing_inst:output_west_empty -> dircc_routing_inst_output_west_bfm:sink_empty
	wire   [0:0] dircc_routing_inst_input_east_bfm_src_valid;          // dircc_routing_inst_input_east_bfm:src_valid -> dircc_routing_inst:input_east_valid
	wire  [31:0] dircc_routing_inst_input_east_bfm_src_data;           // dircc_routing_inst_input_east_bfm:src_data -> dircc_routing_inst:input_east_data
	wire         dircc_routing_inst_input_east_bfm_src_ready;          // dircc_routing_inst:input_east_ready -> dircc_routing_inst_input_east_bfm:src_ready
	wire   [0:0] dircc_routing_inst_input_east_bfm_src_startofpacket;  // dircc_routing_inst_input_east_bfm:src_startofpacket -> dircc_routing_inst:input_east_startofpacket
	wire   [0:0] dircc_routing_inst_input_east_bfm_src_endofpacket;    // dircc_routing_inst_input_east_bfm:src_endofpacket -> dircc_routing_inst:input_east_endofpacket
	wire   [1:0] dircc_routing_inst_input_east_bfm_src_empty;          // dircc_routing_inst_input_east_bfm:src_empty -> dircc_routing_inst:input_east_empty
	wire   [0:0] dircc_routing_inst_input_here_bfm_src_valid;          // dircc_routing_inst_input_here_bfm:src_valid -> dircc_routing_inst:input_here_valid
	wire  [31:0] dircc_routing_inst_input_here_bfm_src_data;           // dircc_routing_inst_input_here_bfm:src_data -> dircc_routing_inst:input_here_data
	wire         dircc_routing_inst_input_here_bfm_src_ready;          // dircc_routing_inst:input_here_ready -> dircc_routing_inst_input_here_bfm:src_ready
	wire   [0:0] dircc_routing_inst_input_here_bfm_src_startofpacket;  // dircc_routing_inst_input_here_bfm:src_startofpacket -> dircc_routing_inst:input_here_startofpacket
	wire   [0:0] dircc_routing_inst_input_here_bfm_src_endofpacket;    // dircc_routing_inst_input_here_bfm:src_endofpacket -> dircc_routing_inst:input_here_endofpacket
	wire   [1:0] dircc_routing_inst_input_here_bfm_src_empty;          // dircc_routing_inst_input_here_bfm:src_empty -> dircc_routing_inst:input_here_empty
	wire   [0:0] dircc_routing_inst_input_north_bfm_src_valid;         // dircc_routing_inst_input_north_bfm:src_valid -> dircc_routing_inst:input_north_valid
	wire  [31:0] dircc_routing_inst_input_north_bfm_src_data;          // dircc_routing_inst_input_north_bfm:src_data -> dircc_routing_inst:input_north_data
	wire         dircc_routing_inst_input_north_bfm_src_ready;         // dircc_routing_inst:input_north_ready -> dircc_routing_inst_input_north_bfm:src_ready
	wire   [0:0] dircc_routing_inst_input_north_bfm_src_startofpacket; // dircc_routing_inst_input_north_bfm:src_startofpacket -> dircc_routing_inst:input_north_startofpacket
	wire   [0:0] dircc_routing_inst_input_north_bfm_src_endofpacket;   // dircc_routing_inst_input_north_bfm:src_endofpacket -> dircc_routing_inst:input_north_endofpacket
	wire   [1:0] dircc_routing_inst_input_north_bfm_src_empty;         // dircc_routing_inst_input_north_bfm:src_empty -> dircc_routing_inst:input_north_empty
	wire   [0:0] dircc_routing_inst_input_south_bfm_src_valid;         // dircc_routing_inst_input_south_bfm:src_valid -> dircc_routing_inst:input_south_valid
	wire  [31:0] dircc_routing_inst_input_south_bfm_src_data;          // dircc_routing_inst_input_south_bfm:src_data -> dircc_routing_inst:input_south_data
	wire         dircc_routing_inst_input_south_bfm_src_ready;         // dircc_routing_inst:input_south_ready -> dircc_routing_inst_input_south_bfm:src_ready
	wire   [0:0] dircc_routing_inst_input_south_bfm_src_startofpacket; // dircc_routing_inst_input_south_bfm:src_startofpacket -> dircc_routing_inst:input_south_startofpacket
	wire   [0:0] dircc_routing_inst_input_south_bfm_src_endofpacket;   // dircc_routing_inst_input_south_bfm:src_endofpacket -> dircc_routing_inst:input_south_endofpacket
	wire   [1:0] dircc_routing_inst_input_south_bfm_src_empty;         // dircc_routing_inst_input_south_bfm:src_empty -> dircc_routing_inst:input_south_empty
	wire   [0:0] dircc_routing_inst_input_west_bfm_src_valid;          // dircc_routing_inst_input_west_bfm:src_valid -> dircc_routing_inst:input_west_valid
	wire  [31:0] dircc_routing_inst_input_west_bfm_src_data;           // dircc_routing_inst_input_west_bfm:src_data -> dircc_routing_inst:input_west_data
	wire         dircc_routing_inst_input_west_bfm_src_ready;          // dircc_routing_inst:input_west_ready -> dircc_routing_inst_input_west_bfm:src_ready
	wire   [0:0] dircc_routing_inst_input_west_bfm_src_startofpacket;  // dircc_routing_inst_input_west_bfm:src_startofpacket -> dircc_routing_inst:input_west_startofpacket
	wire   [0:0] dircc_routing_inst_input_west_bfm_src_endofpacket;    // dircc_routing_inst_input_west_bfm:src_endofpacket -> dircc_routing_inst:input_west_endofpacket
	wire   [1:0] dircc_routing_inst_input_west_bfm_src_empty;          // dircc_routing_inst_input_west_bfm:src_empty -> dircc_routing_inst:input_west_empty
	wire         dircc_routing_inst_clk_bfm_clk_clk;                   // dircc_routing_inst_clk_bfm:clk -> [dircc_routing_inst:clk_clk, dircc_routing_inst_input_east_bfm:clk, dircc_routing_inst_input_here_bfm:clk, dircc_routing_inst_input_north_bfm:clk, dircc_routing_inst_input_south_bfm:clk, dircc_routing_inst_input_west_bfm:clk, dircc_routing_inst_output_east_bfm:clk, dircc_routing_inst_output_here_bfm:clk, dircc_routing_inst_output_north_bfm:clk, dircc_routing_inst_output_south_bfm:clk, dircc_routing_inst_output_west_bfm:clk, dircc_routing_inst_reset_bfm:clk]
	wire  [31:0] dircc_routing_inst_address_bfm_conduit_address;       // dircc_routing_inst_address_bfm:sig_address -> dircc_routing_inst:address_address
	wire         dircc_routing_inst_reset_bfm_reset_reset;             // dircc_routing_inst_reset_bfm:reset -> [dircc_routing_inst:reset_reset_n, dircc_routing_inst_input_east_bfm:reset, dircc_routing_inst_input_here_bfm:reset, dircc_routing_inst_input_north_bfm:reset, dircc_routing_inst_input_south_bfm:reset, dircc_routing_inst_input_west_bfm:reset, dircc_routing_inst_output_east_bfm:reset, dircc_routing_inst_output_here_bfm:reset, dircc_routing_inst_output_north_bfm:reset, dircc_routing_inst_output_south_bfm:reset, dircc_routing_inst_output_west_bfm:reset]

	dircc_routing dircc_routing_inst (
		.address_address            (dircc_routing_inst_address_bfm_conduit_address),       //      address.address
		.clk_clk                    (dircc_routing_inst_clk_bfm_clk_clk),                   //          clk.clk
		.input_east_data            (dircc_routing_inst_input_east_bfm_src_data),           //   input_east.data
		.input_east_valid           (dircc_routing_inst_input_east_bfm_src_valid),          //             .valid
		.input_east_ready           (dircc_routing_inst_input_east_bfm_src_ready),          //             .ready
		.input_east_startofpacket   (dircc_routing_inst_input_east_bfm_src_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (dircc_routing_inst_input_east_bfm_src_endofpacket),    //             .endofpacket
		.input_east_empty           (dircc_routing_inst_input_east_bfm_src_empty),          //             .empty
		.input_here_data            (dircc_routing_inst_input_here_bfm_src_data),           //   input_here.data
		.input_here_valid           (dircc_routing_inst_input_here_bfm_src_valid),          //             .valid
		.input_here_ready           (dircc_routing_inst_input_here_bfm_src_ready),          //             .ready
		.input_here_startofpacket   (dircc_routing_inst_input_here_bfm_src_startofpacket),  //             .startofpacket
		.input_here_endofpacket     (dircc_routing_inst_input_here_bfm_src_endofpacket),    //             .endofpacket
		.input_here_empty           (dircc_routing_inst_input_here_bfm_src_empty),          //             .empty
		.input_north_data           (dircc_routing_inst_input_north_bfm_src_data),          //  input_north.data
		.input_north_valid          (dircc_routing_inst_input_north_bfm_src_valid),         //             .valid
		.input_north_ready          (dircc_routing_inst_input_north_bfm_src_ready),         //             .ready
		.input_north_startofpacket  (dircc_routing_inst_input_north_bfm_src_startofpacket), //             .startofpacket
		.input_north_endofpacket    (dircc_routing_inst_input_north_bfm_src_endofpacket),   //             .endofpacket
		.input_north_empty          (dircc_routing_inst_input_north_bfm_src_empty),         //             .empty
		.input_south_data           (dircc_routing_inst_input_south_bfm_src_data),          //  input_south.data
		.input_south_valid          (dircc_routing_inst_input_south_bfm_src_valid),         //             .valid
		.input_south_ready          (dircc_routing_inst_input_south_bfm_src_ready),         //             .ready
		.input_south_startofpacket  (dircc_routing_inst_input_south_bfm_src_startofpacket), //             .startofpacket
		.input_south_endofpacket    (dircc_routing_inst_input_south_bfm_src_endofpacket),   //             .endofpacket
		.input_south_empty          (dircc_routing_inst_input_south_bfm_src_empty),         //             .empty
		.input_west_data            (dircc_routing_inst_input_west_bfm_src_data),           //   input_west.data
		.input_west_valid           (dircc_routing_inst_input_west_bfm_src_valid),          //             .valid
		.input_west_ready           (dircc_routing_inst_input_west_bfm_src_ready),          //             .ready
		.input_west_startofpacket   (dircc_routing_inst_input_west_bfm_src_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (dircc_routing_inst_input_west_bfm_src_endofpacket),    //             .endofpacket
		.input_west_empty           (dircc_routing_inst_input_west_bfm_src_empty),          //             .empty
		.output_east_data           (dircc_routing_inst_output_east_data),                  //  output_east.data
		.output_east_valid          (dircc_routing_inst_output_east_valid),                 //             .valid
		.output_east_ready          (dircc_routing_inst_output_east_ready),                 //             .ready
		.output_east_startofpacket  (dircc_routing_inst_output_east_startofpacket),         //             .startofpacket
		.output_east_endofpacket    (dircc_routing_inst_output_east_endofpacket),           //             .endofpacket
		.output_east_empty          (dircc_routing_inst_output_east_empty),                 //             .empty
		.output_here_data           (dircc_routing_inst_output_here_data),                  //  output_here.data
		.output_here_valid          (dircc_routing_inst_output_here_valid),                 //             .valid
		.output_here_ready          (dircc_routing_inst_output_here_ready),                 //             .ready
		.output_here_startofpacket  (dircc_routing_inst_output_here_startofpacket),         //             .startofpacket
		.output_here_endofpacket    (dircc_routing_inst_output_here_endofpacket),           //             .endofpacket
		.output_here_empty          (dircc_routing_inst_output_here_empty),                 //             .empty
		.output_north_data          (dircc_routing_inst_output_north_data),                 // output_north.data
		.output_north_valid         (dircc_routing_inst_output_north_valid),                //             .valid
		.output_north_ready         (dircc_routing_inst_output_north_ready),                //             .ready
		.output_north_startofpacket (dircc_routing_inst_output_north_startofpacket),        //             .startofpacket
		.output_north_endofpacket   (dircc_routing_inst_output_north_endofpacket),          //             .endofpacket
		.output_north_empty         (dircc_routing_inst_output_north_empty),                //             .empty
		.output_south_data          (dircc_routing_inst_output_south_data),                 // output_south.data
		.output_south_valid         (dircc_routing_inst_output_south_valid),                //             .valid
		.output_south_ready         (dircc_routing_inst_output_south_ready),                //             .ready
		.output_south_startofpacket (dircc_routing_inst_output_south_startofpacket),        //             .startofpacket
		.output_south_endofpacket   (dircc_routing_inst_output_south_endofpacket),          //             .endofpacket
		.output_south_empty         (dircc_routing_inst_output_south_empty),                //             .empty
		.output_west_data           (dircc_routing_inst_output_west_data),                  //  output_west.data
		.output_west_valid          (dircc_routing_inst_output_west_valid),                 //             .valid
		.output_west_ready          (dircc_routing_inst_output_west_ready),                 //             .ready
		.output_west_startofpacket  (dircc_routing_inst_output_west_startofpacket),         //             .startofpacket
		.output_west_endofpacket    (dircc_routing_inst_output_west_endofpacket),           //             .endofpacket
		.output_west_empty          (dircc_routing_inst_output_west_empty),                 //             .empty
		.reset_reset_n              (dircc_routing_inst_reset_bfm_reset_reset)              //        reset.reset_n
	);

	altera_conduit_bfm dircc_routing_inst_address_bfm (
		.sig_address (dircc_routing_inst_address_bfm_conduit_address)  // conduit.address
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dircc_routing_inst_clk_bfm (
		.clk (dircc_routing_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dircc_routing_inst_input_east_bfm (
		.clk               (dircc_routing_inst_clk_bfm_clk_clk),                  //       clk.clk
		.reset             (~dircc_routing_inst_reset_bfm_reset_reset),           // clk_reset.reset
		.src_data          (dircc_routing_inst_input_east_bfm_src_data),          //       src.data
		.src_valid         (dircc_routing_inst_input_east_bfm_src_valid),         //          .valid
		.src_ready         (dircc_routing_inst_input_east_bfm_src_ready),         //          .ready
		.src_startofpacket (dircc_routing_inst_input_east_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (dircc_routing_inst_input_east_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (dircc_routing_inst_input_east_bfm_src_empty),         //          .empty
		.src_channel       (),                                                    // (terminated)
		.src_error         ()                                                     // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (1)
	) dircc_routing_inst_input_here_bfm (
		.clk               (dircc_routing_inst_clk_bfm_clk_clk),                  //       clk.clk
		.reset             (~dircc_routing_inst_reset_bfm_reset_reset),           // clk_reset.reset
		.src_data          (dircc_routing_inst_input_here_bfm_src_data),          //       src.data
		.src_valid         (dircc_routing_inst_input_here_bfm_src_valid),         //          .valid
		.src_ready         (dircc_routing_inst_input_here_bfm_src_ready),         //          .ready
		.src_startofpacket (dircc_routing_inst_input_here_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (dircc_routing_inst_input_here_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (dircc_routing_inst_input_here_bfm_src_empty),         //          .empty
		.src_channel       (),                                                    // (terminated)
		.src_error         ()                                                     // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (2)
	) dircc_routing_inst_input_north_bfm (
		.clk               (dircc_routing_inst_clk_bfm_clk_clk),                   //       clk.clk
		.reset             (~dircc_routing_inst_reset_bfm_reset_reset),            // clk_reset.reset
		.src_data          (dircc_routing_inst_input_north_bfm_src_data),          //       src.data
		.src_valid         (dircc_routing_inst_input_north_bfm_src_valid),         //          .valid
		.src_ready         (dircc_routing_inst_input_north_bfm_src_ready),         //          .ready
		.src_startofpacket (dircc_routing_inst_input_north_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (dircc_routing_inst_input_north_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (dircc_routing_inst_input_north_bfm_src_empty),         //          .empty
		.src_channel       (),                                                     // (terminated)
		.src_error         ()                                                      // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (3)
	) dircc_routing_inst_input_south_bfm (
		.clk               (dircc_routing_inst_clk_bfm_clk_clk),                   //       clk.clk
		.reset             (~dircc_routing_inst_reset_bfm_reset_reset),            // clk_reset.reset
		.src_data          (dircc_routing_inst_input_south_bfm_src_data),          //       src.data
		.src_valid         (dircc_routing_inst_input_south_bfm_src_valid),         //          .valid
		.src_ready         (dircc_routing_inst_input_south_bfm_src_ready),         //          .ready
		.src_startofpacket (dircc_routing_inst_input_south_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (dircc_routing_inst_input_south_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (dircc_routing_inst_input_south_bfm_src_empty),         //          .empty
		.src_channel       (),                                                     // (terminated)
		.src_error         ()                                                      // (terminated)
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (4)
	) dircc_routing_inst_input_west_bfm (
		.clk               (dircc_routing_inst_clk_bfm_clk_clk),                  //       clk.clk
		.reset             (~dircc_routing_inst_reset_bfm_reset_reset),           // clk_reset.reset
		.src_data          (dircc_routing_inst_input_west_bfm_src_data),          //       src.data
		.src_valid         (dircc_routing_inst_input_west_bfm_src_valid),         //          .valid
		.src_ready         (dircc_routing_inst_input_west_bfm_src_ready),         //          .ready
		.src_startofpacket (dircc_routing_inst_input_west_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (dircc_routing_inst_input_west_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (dircc_routing_inst_input_west_bfm_src_empty),         //          .empty
		.src_channel       (),                                                    // (terminated)
		.src_error         ()                                                     // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dircc_routing_inst_output_east_bfm (
		.clk                (dircc_routing_inst_clk_bfm_clk_clk),           //       clk.clk
		.reset              (~dircc_routing_inst_reset_bfm_reset_reset),    // clk_reset.reset
		.sink_data          (dircc_routing_inst_output_east_data),          //      sink.data
		.sink_valid         (dircc_routing_inst_output_east_valid),         //          .valid
		.sink_ready         (dircc_routing_inst_output_east_ready),         //          .ready
		.sink_startofpacket (dircc_routing_inst_output_east_startofpacket), //          .startofpacket
		.sink_endofpacket   (dircc_routing_inst_output_east_endofpacket),   //          .endofpacket
		.sink_empty         (dircc_routing_inst_output_east_empty),         //          .empty
		.sink_channel       (1'b0),                                         // (terminated)
		.sink_error         (1'b0)                                          // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (1)
	) dircc_routing_inst_output_here_bfm (
		.clk                (dircc_routing_inst_clk_bfm_clk_clk),           //       clk.clk
		.reset              (~dircc_routing_inst_reset_bfm_reset_reset),    // clk_reset.reset
		.sink_data          (dircc_routing_inst_output_here_data),          //      sink.data
		.sink_valid         (dircc_routing_inst_output_here_valid),         //          .valid
		.sink_ready         (dircc_routing_inst_output_here_ready),         //          .ready
		.sink_startofpacket (dircc_routing_inst_output_here_startofpacket), //          .startofpacket
		.sink_endofpacket   (dircc_routing_inst_output_here_endofpacket),   //          .endofpacket
		.sink_empty         (dircc_routing_inst_output_here_empty),         //          .empty
		.sink_channel       (1'b0),                                         // (terminated)
		.sink_error         (1'b0)                                          // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (2)
	) dircc_routing_inst_output_north_bfm (
		.clk                (dircc_routing_inst_clk_bfm_clk_clk),            //       clk.clk
		.reset              (~dircc_routing_inst_reset_bfm_reset_reset),     // clk_reset.reset
		.sink_data          (dircc_routing_inst_output_north_data),          //      sink.data
		.sink_valid         (dircc_routing_inst_output_north_valid),         //          .valid
		.sink_ready         (dircc_routing_inst_output_north_ready),         //          .ready
		.sink_startofpacket (dircc_routing_inst_output_north_startofpacket), //          .startofpacket
		.sink_endofpacket   (dircc_routing_inst_output_north_endofpacket),   //          .endofpacket
		.sink_empty         (dircc_routing_inst_output_north_empty),         //          .empty
		.sink_channel       (1'b0),                                          // (terminated)
		.sink_error         (1'b0)                                           // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (3)
	) dircc_routing_inst_output_south_bfm (
		.clk                (dircc_routing_inst_clk_bfm_clk_clk),            //       clk.clk
		.reset              (~dircc_routing_inst_reset_bfm_reset_reset),     // clk_reset.reset
		.sink_data          (dircc_routing_inst_output_south_data),          //      sink.data
		.sink_valid         (dircc_routing_inst_output_south_valid),         //          .valid
		.sink_ready         (dircc_routing_inst_output_south_ready),         //          .ready
		.sink_startofpacket (dircc_routing_inst_output_south_startofpacket), //          .startofpacket
		.sink_endofpacket   (dircc_routing_inst_output_south_endofpacket),   //          .endofpacket
		.sink_empty         (dircc_routing_inst_output_south_empty),         //          .empty
		.sink_channel       (1'b0),                                          // (terminated)
		.sink_error         (1'b0)                                           // (terminated)
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (4)
	) dircc_routing_inst_output_west_bfm (
		.clk                (dircc_routing_inst_clk_bfm_clk_clk),           //       clk.clk
		.reset              (~dircc_routing_inst_reset_bfm_reset_reset),    // clk_reset.reset
		.sink_data          (dircc_routing_inst_output_west_data),          //      sink.data
		.sink_valid         (dircc_routing_inst_output_west_valid),         //          .valid
		.sink_ready         (dircc_routing_inst_output_west_ready),         //          .ready
		.sink_startofpacket (dircc_routing_inst_output_west_startofpacket), //          .startofpacket
		.sink_endofpacket   (dircc_routing_inst_output_west_endofpacket),   //          .endofpacket
		.sink_empty         (dircc_routing_inst_output_west_empty),         //          .empty
		.sink_channel       (1'b0),                                         // (terminated)
		.sink_error         (1'b0)                                          // (terminated)
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dircc_routing_inst_reset_bfm (
		.reset (dircc_routing_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dircc_routing_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
