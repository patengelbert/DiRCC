// dircc_processing_counter_test_sys.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_processing_counter_test_sys (
		input  wire        clk_clk,                  //            clk.clk
		output wire [15:0] east_0_mem_readdata,      //     east_0_mem.readdata
		input  wire [1:0]  east_0_mem_address,       //               .address
		input  wire        east_0_mem_read_n,        //               .read_n
		output wire [15:0] east_1_mem_readdata,      //     east_1_mem.readdata
		input  wire [1:0]  east_1_mem_address,       //               .address
		input  wire        east_1_mem_read_n,        //               .read_n
		input  wire [14:0] node_0_mem_address,       //     node_0_mem.address
		output wire [15:0] node_0_mem_readdata,      //               .readdata
		input  wire        node_0_mem_write,         //               .write
		input  wire [15:0] node_0_mem_writedata,     //               .writedata
		input  wire [14:0] node_1_mem_address,       //     node_1_mem.address
		output wire [15:0] node_1_mem_readdata,      //               .readdata
		input  wire        node_1_mem_write,         //               .write
		input  wire [15:0] node_1_mem_writedata,     //               .writedata
		input  wire [14:0] node_65536_mem_address,   // node_65536_mem.address
		output wire [15:0] node_65536_mem_readdata,  //               .readdata
		input  wire        node_65536_mem_write,     //               .write
		input  wire [15:0] node_65536_mem_writedata, //               .writedata
		input  wire [14:0] node_65537_mem_address,   // node_65537_mem.address
		output wire [15:0] node_65537_mem_readdata,  //               .readdata
		input  wire        node_65537_mem_write,     //               .write
		input  wire [15:0] node_65537_mem_writedata, //               .writedata
		output wire [15:0] north_0_mem_readdata,     //    north_0_mem.readdata
		input  wire [1:0]  north_0_mem_address,      //               .address
		input  wire        north_0_mem_read_n,       //               .read_n
		output wire [15:0] north_1_mem_readdata,     //    north_1_mem.readdata
		input  wire [1:0]  north_1_mem_address,      //               .address
		input  wire        north_1_mem_read_n,       //               .read_n
		input  wire        reset_reset_n,            //          reset.reset_n
		output wire [15:0] south_0_mem_readdata,     //    south_0_mem.readdata
		input  wire [1:0]  south_0_mem_address,      //               .address
		input  wire        south_0_mem_read_n,       //               .read_n
		output wire [15:0] south_1_mem_readdata,     //    south_1_mem.readdata
		input  wire [1:0]  south_1_mem_address,      //               .address
		input  wire        south_1_mem_read_n,       //               .read_n
		output wire [15:0] west_0_mem_readdata,      //     west_0_mem.readdata
		input  wire [1:0]  west_0_mem_address,       //               .address
		input  wire        west_0_mem_read_n,        //               .read_n
		output wire [15:0] west_1_mem_readdata,      //     west_1_mem.readdata
		input  wire [1:0]  west_1_mem_address,       //               .address
		input  wire        west_1_mem_read_n         //               .read_n
	);

	wire         node_0_output_east_valid;              // node_0:output_east_valid -> node_1:input_west_valid
	wire  [31:0] node_0_output_east_data;               // node_0:output_east_data -> node_1:input_west_data
	wire         node_0_output_east_ready;              // node_1:input_west_ready -> node_0:output_east_ready
	wire         node_0_output_east_startofpacket;      // node_0:output_east_startofpacket -> node_1:input_west_startofpacket
	wire         node_0_output_east_endofpacket;        // node_0:output_east_endofpacket -> node_1:input_west_endofpacket
	wire   [1:0] node_0_output_east_empty;              // node_0:output_east_empty -> node_1:input_west_empty
	wire         node_65536_output_east_valid;          // node_65536:output_east_valid -> node_65537:input_west_valid
	wire  [31:0] node_65536_output_east_data;           // node_65536:output_east_data -> node_65537:input_west_data
	wire         node_65536_output_east_ready;          // node_65537:input_west_ready -> node_65536:output_east_ready
	wire         node_65536_output_east_startofpacket;  // node_65536:output_east_startofpacket -> node_65537:input_west_startofpacket
	wire         node_65536_output_east_endofpacket;    // node_65536:output_east_endofpacket -> node_65537:input_west_endofpacket
	wire   [1:0] node_65536_output_east_empty;          // node_65536:output_east_empty -> node_65537:input_west_empty
	wire         node_1_output_east_valid;              // node_1:output_east_valid -> terminal_east_0:valid
	wire  [31:0] node_1_output_east_data;               // node_1:output_east_data -> terminal_east_0:data
	wire         node_1_output_east_ready;              // terminal_east_0:ready -> node_1:output_east_ready
	wire         node_1_output_east_startofpacket;      // node_1:output_east_startofpacket -> terminal_east_0:startofpacket
	wire         node_1_output_east_endofpacket;        // node_1:output_east_endofpacket -> terminal_east_0:endofpacket
	wire   [1:0] node_1_output_east_empty;              // node_1:output_east_empty -> terminal_east_0:empty
	wire         node_65537_output_east_valid;          // node_65537:output_east_valid -> terminal_east_1:valid
	wire  [31:0] node_65537_output_east_data;           // node_65537:output_east_data -> terminal_east_1:data
	wire         node_65537_output_east_ready;          // terminal_east_1:ready -> node_65537:output_east_ready
	wire         node_65537_output_east_startofpacket;  // node_65537:output_east_startofpacket -> terminal_east_1:startofpacket
	wire         node_65537_output_east_endofpacket;    // node_65537:output_east_endofpacket -> terminal_east_1:endofpacket
	wire   [1:0] node_65537_output_east_empty;          // node_65537:output_east_empty -> terminal_east_1:empty
	wire         node_65537_output_north_valid;         // node_65537:output_north_valid -> node_1:input_south_valid
	wire  [31:0] node_65537_output_north_data;          // node_65537:output_north_data -> node_1:input_south_data
	wire         node_65537_output_north_ready;         // node_1:input_south_ready -> node_65537:output_north_ready
	wire         node_65537_output_north_startofpacket; // node_65537:output_north_startofpacket -> node_1:input_south_startofpacket
	wire         node_65537_output_north_endofpacket;   // node_65537:output_north_endofpacket -> node_1:input_south_endofpacket
	wire   [1:0] node_65537_output_north_empty;         // node_65537:output_north_empty -> node_1:input_south_empty
	wire         node_65536_output_north_valid;         // node_65536:output_north_valid -> node_0:input_south_valid
	wire  [31:0] node_65536_output_north_data;          // node_65536:output_north_data -> node_0:input_south_data
	wire         node_65536_output_north_ready;         // node_0:input_south_ready -> node_65536:output_north_ready
	wire         node_65536_output_north_startofpacket; // node_65536:output_north_startofpacket -> node_0:input_south_startofpacket
	wire         node_65536_output_north_endofpacket;   // node_65536:output_north_endofpacket -> node_0:input_south_endofpacket
	wire   [1:0] node_65536_output_north_empty;         // node_65536:output_north_empty -> node_0:input_south_empty
	wire         node_0_output_north_valid;             // node_0:output_north_valid -> terminal_north_0:valid
	wire  [31:0] node_0_output_north_data;              // node_0:output_north_data -> terminal_north_0:data
	wire         node_0_output_north_ready;             // terminal_north_0:ready -> node_0:output_north_ready
	wire         node_0_output_north_startofpacket;     // node_0:output_north_startofpacket -> terminal_north_0:startofpacket
	wire         node_0_output_north_endofpacket;       // node_0:output_north_endofpacket -> terminal_north_0:endofpacket
	wire   [1:0] node_0_output_north_empty;             // node_0:output_north_empty -> terminal_north_0:empty
	wire         node_1_output_north_valid;             // node_1:output_north_valid -> terminal_north_1:valid
	wire  [31:0] node_1_output_north_data;              // node_1:output_north_data -> terminal_north_1:data
	wire         node_1_output_north_ready;             // terminal_north_1:ready -> node_1:output_north_ready
	wire         node_1_output_north_startofpacket;     // node_1:output_north_startofpacket -> terminal_north_1:startofpacket
	wire         node_1_output_north_endofpacket;       // node_1:output_north_endofpacket -> terminal_north_1:endofpacket
	wire   [1:0] node_1_output_north_empty;             // node_1:output_north_empty -> terminal_north_1:empty
	wire         node_1_output_south_valid;             // node_1:output_south_valid -> node_65537:input_north_valid
	wire  [31:0] node_1_output_south_data;              // node_1:output_south_data -> node_65537:input_north_data
	wire         node_1_output_south_ready;             // node_65537:input_north_ready -> node_1:output_south_ready
	wire         node_1_output_south_startofpacket;     // node_1:output_south_startofpacket -> node_65537:input_north_startofpacket
	wire         node_1_output_south_endofpacket;       // node_1:output_south_endofpacket -> node_65537:input_north_endofpacket
	wire   [1:0] node_1_output_south_empty;             // node_1:output_south_empty -> node_65537:input_north_empty
	wire         node_0_output_south_valid;             // node_0:output_south_valid -> node_65536:input_north_valid
	wire  [31:0] node_0_output_south_data;              // node_0:output_south_data -> node_65536:input_north_data
	wire         node_0_output_south_ready;             // node_65536:input_north_ready -> node_0:output_south_ready
	wire         node_0_output_south_startofpacket;     // node_0:output_south_startofpacket -> node_65536:input_north_startofpacket
	wire         node_0_output_south_endofpacket;       // node_0:output_south_endofpacket -> node_65536:input_north_endofpacket
	wire   [1:0] node_0_output_south_empty;             // node_0:output_south_empty -> node_65536:input_north_empty
	wire         node_65536_output_south_valid;         // node_65536:output_south_valid -> terminal_south_0:valid
	wire  [31:0] node_65536_output_south_data;          // node_65536:output_south_data -> terminal_south_0:data
	wire         node_65536_output_south_ready;         // terminal_south_0:ready -> node_65536:output_south_ready
	wire         node_65536_output_south_startofpacket; // node_65536:output_south_startofpacket -> terminal_south_0:startofpacket
	wire         node_65536_output_south_endofpacket;   // node_65536:output_south_endofpacket -> terminal_south_0:endofpacket
	wire   [1:0] node_65536_output_south_empty;         // node_65536:output_south_empty -> terminal_south_0:empty
	wire         node_65537_output_south_valid;         // node_65537:output_south_valid -> terminal_south_1:valid
	wire  [31:0] node_65537_output_south_data;          // node_65537:output_south_data -> terminal_south_1:data
	wire         node_65537_output_south_ready;         // terminal_south_1:ready -> node_65537:output_south_ready
	wire         node_65537_output_south_startofpacket; // node_65537:output_south_startofpacket -> terminal_south_1:startofpacket
	wire         node_65537_output_south_endofpacket;   // node_65537:output_south_endofpacket -> terminal_south_1:endofpacket
	wire   [1:0] node_65537_output_south_empty;         // node_65537:output_south_empty -> terminal_south_1:empty
	wire         node_1_output_west_valid;              // node_1:output_west_valid -> node_0:input_east_valid
	wire  [31:0] node_1_output_west_data;               // node_1:output_west_data -> node_0:input_east_data
	wire         node_1_output_west_ready;              // node_0:input_east_ready -> node_1:output_west_ready
	wire         node_1_output_west_startofpacket;      // node_1:output_west_startofpacket -> node_0:input_east_startofpacket
	wire         node_1_output_west_endofpacket;        // node_1:output_west_endofpacket -> node_0:input_east_endofpacket
	wire   [1:0] node_1_output_west_empty;              // node_1:output_west_empty -> node_0:input_east_empty
	wire         node_65537_output_west_valid;          // node_65537:output_west_valid -> node_65536:input_east_valid
	wire  [31:0] node_65537_output_west_data;           // node_65537:output_west_data -> node_65536:input_east_data
	wire         node_65537_output_west_ready;          // node_65536:input_east_ready -> node_65537:output_west_ready
	wire         node_65537_output_west_startofpacket;  // node_65537:output_west_startofpacket -> node_65536:input_east_startofpacket
	wire         node_65537_output_west_endofpacket;    // node_65537:output_west_endofpacket -> node_65536:input_east_endofpacket
	wire   [1:0] node_65537_output_west_empty;          // node_65537:output_west_empty -> node_65536:input_east_empty
	wire         node_0_output_west_valid;              // node_0:output_west_valid -> terminal_west_0:valid
	wire  [31:0] node_0_output_west_data;               // node_0:output_west_data -> terminal_west_0:data
	wire         node_0_output_west_ready;              // terminal_west_0:ready -> node_0:output_west_ready
	wire         node_0_output_west_startofpacket;      // node_0:output_west_startofpacket -> terminal_west_0:startofpacket
	wire         node_0_output_west_endofpacket;        // node_0:output_west_endofpacket -> terminal_west_0:endofpacket
	wire   [1:0] node_0_output_west_empty;              // node_0:output_west_empty -> terminal_west_0:empty
	wire         node_65536_output_west_valid;          // node_65536:output_west_valid -> terminal_west_1:valid
	wire  [31:0] node_65536_output_west_data;           // node_65536:output_west_data -> terminal_west_1:data
	wire         node_65536_output_west_ready;          // terminal_west_1:ready -> node_65536:output_west_ready
	wire         node_65536_output_west_startofpacket;  // node_65536:output_west_startofpacket -> terminal_west_1:startofpacket
	wire         node_65536_output_west_endofpacket;    // node_65536:output_west_endofpacket -> terminal_west_1:endofpacket
	wire   [1:0] node_65536_output_west_empty;          // node_65536:output_west_empty -> terminal_west_1:empty
	wire         rst_controller_reset_out_reset;        // rst_controller:reset_out -> [terminal_east_0:reset_n, terminal_east_1:reset_n, terminal_north_0:reset_n, terminal_north_1:reset_n, terminal_south_0:reset_n, terminal_south_1:reset_n, terminal_west_0:reset_n, terminal_west_1:reset_n]

	dircc_processing_counter_test_sys_node_0 node_0 (
		.clk_clk                    (clk_clk),                               //            clk.clk
		.input_east_data            (node_1_output_west_data),               //     input_east.data
		.input_east_valid           (node_1_output_west_valid),              //               .valid
		.input_east_ready           (node_1_output_west_ready),              //               .ready
		.input_east_startofpacket   (node_1_output_west_startofpacket),      //               .startofpacket
		.input_east_endofpacket     (node_1_output_west_endofpacket),        //               .endofpacket
		.input_east_empty           (node_1_output_west_empty),              //               .empty
		.input_north_data           (),                                      //    input_north.data
		.input_north_valid          (),                                      //               .valid
		.input_north_ready          (),                                      //               .ready
		.input_north_startofpacket  (),                                      //               .startofpacket
		.input_north_endofpacket    (),                                      //               .endofpacket
		.input_north_empty          (),                                      //               .empty
		.input_south_data           (node_65536_output_north_data),          //    input_south.data
		.input_south_valid          (node_65536_output_north_valid),         //               .valid
		.input_south_ready          (node_65536_output_north_ready),         //               .ready
		.input_south_startofpacket  (node_65536_output_north_startofpacket), //               .startofpacket
		.input_south_endofpacket    (node_65536_output_north_endofpacket),   //               .endofpacket
		.input_south_empty          (node_65536_output_north_empty),         //               .empty
		.input_west_data            (),                                      //     input_west.data
		.input_west_valid           (),                                      //               .valid
		.input_west_ready           (),                                      //               .ready
		.input_west_startofpacket   (),                                      //               .startofpacket
		.input_west_endofpacket     (),                                      //               .endofpacket
		.input_west_empty           (),                                      //               .empty
		.output_east_data           (node_0_output_east_data),               //    output_east.data
		.output_east_valid          (node_0_output_east_valid),              //               .valid
		.output_east_ready          (node_0_output_east_ready),              //               .ready
		.output_east_startofpacket  (node_0_output_east_startofpacket),      //               .startofpacket
		.output_east_endofpacket    (node_0_output_east_endofpacket),        //               .endofpacket
		.output_east_empty          (node_0_output_east_empty),              //               .empty
		.output_north_data          (node_0_output_north_data),              //   output_north.data
		.output_north_valid         (node_0_output_north_valid),             //               .valid
		.output_north_ready         (node_0_output_north_ready),             //               .ready
		.output_north_startofpacket (node_0_output_north_startofpacket),     //               .startofpacket
		.output_north_endofpacket   (node_0_output_north_endofpacket),       //               .endofpacket
		.output_north_empty         (node_0_output_north_empty),             //               .empty
		.output_south_data          (node_0_output_south_data),              //   output_south.data
		.output_south_valid         (node_0_output_south_valid),             //               .valid
		.output_south_ready         (node_0_output_south_ready),             //               .ready
		.output_south_startofpacket (node_0_output_south_startofpacket),     //               .startofpacket
		.output_south_endofpacket   (node_0_output_south_endofpacket),       //               .endofpacket
		.output_south_empty         (node_0_output_south_empty),             //               .empty
		.output_west_data           (node_0_output_west_data),               //    output_west.data
		.output_west_valid          (node_0_output_west_valid),              //               .valid
		.output_west_ready          (node_0_output_west_ready),              //               .ready
		.output_west_startofpacket  (node_0_output_west_startofpacket),      //               .startofpacket
		.output_west_endofpacket    (node_0_output_west_endofpacket),        //               .endofpacket
		.output_west_empty          (node_0_output_west_empty),              //               .empty
		.processing_mem_address     (node_0_mem_address),                    // processing_mem.address
		.processing_mem_readdata    (node_0_mem_readdata),                   //               .readdata
		.processing_mem_write       (node_0_mem_write),                      //               .write
		.processing_mem_writedata   (node_0_mem_writedata),                  //               .writedata
		.reset_reset_n              (reset_reset_n)                          //          reset.reset_n
	);

	dircc_processing_counter_test_sys_node_1 node_1 (
		.clk_clk                    (clk_clk),                               //            clk.clk
		.input_east_data            (),                                      //     input_east.data
		.input_east_valid           (),                                      //               .valid
		.input_east_ready           (),                                      //               .ready
		.input_east_startofpacket   (),                                      //               .startofpacket
		.input_east_endofpacket     (),                                      //               .endofpacket
		.input_east_empty           (),                                      //               .empty
		.input_north_data           (),                                      //    input_north.data
		.input_north_valid          (),                                      //               .valid
		.input_north_ready          (),                                      //               .ready
		.input_north_startofpacket  (),                                      //               .startofpacket
		.input_north_endofpacket    (),                                      //               .endofpacket
		.input_north_empty          (),                                      //               .empty
		.input_south_data           (node_65537_output_north_data),          //    input_south.data
		.input_south_valid          (node_65537_output_north_valid),         //               .valid
		.input_south_ready          (node_65537_output_north_ready),         //               .ready
		.input_south_startofpacket  (node_65537_output_north_startofpacket), //               .startofpacket
		.input_south_endofpacket    (node_65537_output_north_endofpacket),   //               .endofpacket
		.input_south_empty          (node_65537_output_north_empty),         //               .empty
		.input_west_data            (node_0_output_east_data),               //     input_west.data
		.input_west_valid           (node_0_output_east_valid),              //               .valid
		.input_west_ready           (node_0_output_east_ready),              //               .ready
		.input_west_startofpacket   (node_0_output_east_startofpacket),      //               .startofpacket
		.input_west_endofpacket     (node_0_output_east_endofpacket),        //               .endofpacket
		.input_west_empty           (node_0_output_east_empty),              //               .empty
		.output_east_data           (node_1_output_east_data),               //    output_east.data
		.output_east_valid          (node_1_output_east_valid),              //               .valid
		.output_east_ready          (node_1_output_east_ready),              //               .ready
		.output_east_startofpacket  (node_1_output_east_startofpacket),      //               .startofpacket
		.output_east_endofpacket    (node_1_output_east_endofpacket),        //               .endofpacket
		.output_east_empty          (node_1_output_east_empty),              //               .empty
		.output_north_data          (node_1_output_north_data),              //   output_north.data
		.output_north_valid         (node_1_output_north_valid),             //               .valid
		.output_north_ready         (node_1_output_north_ready),             //               .ready
		.output_north_startofpacket (node_1_output_north_startofpacket),     //               .startofpacket
		.output_north_endofpacket   (node_1_output_north_endofpacket),       //               .endofpacket
		.output_north_empty         (node_1_output_north_empty),             //               .empty
		.output_south_data          (node_1_output_south_data),              //   output_south.data
		.output_south_valid         (node_1_output_south_valid),             //               .valid
		.output_south_ready         (node_1_output_south_ready),             //               .ready
		.output_south_startofpacket (node_1_output_south_startofpacket),     //               .startofpacket
		.output_south_endofpacket   (node_1_output_south_endofpacket),       //               .endofpacket
		.output_south_empty         (node_1_output_south_empty),             //               .empty
		.output_west_data           (node_1_output_west_data),               //    output_west.data
		.output_west_valid          (node_1_output_west_valid),              //               .valid
		.output_west_ready          (node_1_output_west_ready),              //               .ready
		.output_west_startofpacket  (node_1_output_west_startofpacket),      //               .startofpacket
		.output_west_endofpacket    (node_1_output_west_endofpacket),        //               .endofpacket
		.output_west_empty          (node_1_output_west_empty),              //               .empty
		.processing_mem_address     (node_1_mem_address),                    // processing_mem.address
		.processing_mem_readdata    (node_1_mem_readdata),                   //               .readdata
		.processing_mem_write       (node_1_mem_write),                      //               .write
		.processing_mem_writedata   (node_1_mem_writedata),                  //               .writedata
		.reset_reset_n              (reset_reset_n)                          //          reset.reset_n
	);

	dircc_processing_counter_test_sys_node_65536 node_65536 (
		.clk_clk                    (clk_clk),                               //            clk.clk
		.input_east_data            (node_65537_output_west_data),           //     input_east.data
		.input_east_valid           (node_65537_output_west_valid),          //               .valid
		.input_east_ready           (node_65537_output_west_ready),          //               .ready
		.input_east_startofpacket   (node_65537_output_west_startofpacket),  //               .startofpacket
		.input_east_endofpacket     (node_65537_output_west_endofpacket),    //               .endofpacket
		.input_east_empty           (node_65537_output_west_empty),          //               .empty
		.input_north_data           (node_0_output_south_data),              //    input_north.data
		.input_north_valid          (node_0_output_south_valid),             //               .valid
		.input_north_ready          (node_0_output_south_ready),             //               .ready
		.input_north_startofpacket  (node_0_output_south_startofpacket),     //               .startofpacket
		.input_north_endofpacket    (node_0_output_south_endofpacket),       //               .endofpacket
		.input_north_empty          (node_0_output_south_empty),             //               .empty
		.input_south_data           (),                                      //    input_south.data
		.input_south_valid          (),                                      //               .valid
		.input_south_ready          (),                                      //               .ready
		.input_south_startofpacket  (),                                      //               .startofpacket
		.input_south_endofpacket    (),                                      //               .endofpacket
		.input_south_empty          (),                                      //               .empty
		.input_west_data            (),                                      //     input_west.data
		.input_west_valid           (),                                      //               .valid
		.input_west_ready           (),                                      //               .ready
		.input_west_startofpacket   (),                                      //               .startofpacket
		.input_west_endofpacket     (),                                      //               .endofpacket
		.input_west_empty           (),                                      //               .empty
		.output_east_data           (node_65536_output_east_data),           //    output_east.data
		.output_east_valid          (node_65536_output_east_valid),          //               .valid
		.output_east_ready          (node_65536_output_east_ready),          //               .ready
		.output_east_startofpacket  (node_65536_output_east_startofpacket),  //               .startofpacket
		.output_east_endofpacket    (node_65536_output_east_endofpacket),    //               .endofpacket
		.output_east_empty          (node_65536_output_east_empty),          //               .empty
		.output_north_data          (node_65536_output_north_data),          //   output_north.data
		.output_north_valid         (node_65536_output_north_valid),         //               .valid
		.output_north_ready         (node_65536_output_north_ready),         //               .ready
		.output_north_startofpacket (node_65536_output_north_startofpacket), //               .startofpacket
		.output_north_endofpacket   (node_65536_output_north_endofpacket),   //               .endofpacket
		.output_north_empty         (node_65536_output_north_empty),         //               .empty
		.output_south_data          (node_65536_output_south_data),          //   output_south.data
		.output_south_valid         (node_65536_output_south_valid),         //               .valid
		.output_south_ready         (node_65536_output_south_ready),         //               .ready
		.output_south_startofpacket (node_65536_output_south_startofpacket), //               .startofpacket
		.output_south_endofpacket   (node_65536_output_south_endofpacket),   //               .endofpacket
		.output_south_empty         (node_65536_output_south_empty),         //               .empty
		.output_west_data           (node_65536_output_west_data),           //    output_west.data
		.output_west_valid          (node_65536_output_west_valid),          //               .valid
		.output_west_ready          (node_65536_output_west_ready),          //               .ready
		.output_west_startofpacket  (node_65536_output_west_startofpacket),  //               .startofpacket
		.output_west_endofpacket    (node_65536_output_west_endofpacket),    //               .endofpacket
		.output_west_empty          (node_65536_output_west_empty),          //               .empty
		.processing_mem_address     (node_65536_mem_address),                // processing_mem.address
		.processing_mem_readdata    (node_65536_mem_readdata),               //               .readdata
		.processing_mem_write       (node_65536_mem_write),                  //               .write
		.processing_mem_writedata   (node_65536_mem_writedata),              //               .writedata
		.reset_reset_n              (reset_reset_n)                          //          reset.reset_n
	);

	dircc_processing_counter_test_sys_node_65537 node_65537 (
		.clk_clk                    (clk_clk),                               //            clk.clk
		.input_east_data            (),                                      //     input_east.data
		.input_east_valid           (),                                      //               .valid
		.input_east_ready           (),                                      //               .ready
		.input_east_startofpacket   (),                                      //               .startofpacket
		.input_east_endofpacket     (),                                      //               .endofpacket
		.input_east_empty           (),                                      //               .empty
		.input_north_data           (node_1_output_south_data),              //    input_north.data
		.input_north_valid          (node_1_output_south_valid),             //               .valid
		.input_north_ready          (node_1_output_south_ready),             //               .ready
		.input_north_startofpacket  (node_1_output_south_startofpacket),     //               .startofpacket
		.input_north_endofpacket    (node_1_output_south_endofpacket),       //               .endofpacket
		.input_north_empty          (node_1_output_south_empty),             //               .empty
		.input_south_data           (),                                      //    input_south.data
		.input_south_valid          (),                                      //               .valid
		.input_south_ready          (),                                      //               .ready
		.input_south_startofpacket  (),                                      //               .startofpacket
		.input_south_endofpacket    (),                                      //               .endofpacket
		.input_south_empty          (),                                      //               .empty
		.input_west_data            (node_65536_output_east_data),           //     input_west.data
		.input_west_valid           (node_65536_output_east_valid),          //               .valid
		.input_west_ready           (node_65536_output_east_ready),          //               .ready
		.input_west_startofpacket   (node_65536_output_east_startofpacket),  //               .startofpacket
		.input_west_endofpacket     (node_65536_output_east_endofpacket),    //               .endofpacket
		.input_west_empty           (node_65536_output_east_empty),          //               .empty
		.output_east_data           (node_65537_output_east_data),           //    output_east.data
		.output_east_valid          (node_65537_output_east_valid),          //               .valid
		.output_east_ready          (node_65537_output_east_ready),          //               .ready
		.output_east_startofpacket  (node_65537_output_east_startofpacket),  //               .startofpacket
		.output_east_endofpacket    (node_65537_output_east_endofpacket),    //               .endofpacket
		.output_east_empty          (node_65537_output_east_empty),          //               .empty
		.output_north_data          (node_65537_output_north_data),          //   output_north.data
		.output_north_valid         (node_65537_output_north_valid),         //               .valid
		.output_north_ready         (node_65537_output_north_ready),         //               .ready
		.output_north_startofpacket (node_65537_output_north_startofpacket), //               .startofpacket
		.output_north_endofpacket   (node_65537_output_north_endofpacket),   //               .endofpacket
		.output_north_empty         (node_65537_output_north_empty),         //               .empty
		.output_south_data          (node_65537_output_south_data),          //   output_south.data
		.output_south_valid         (node_65537_output_south_valid),         //               .valid
		.output_south_ready         (node_65537_output_south_ready),         //               .ready
		.output_south_startofpacket (node_65537_output_south_startofpacket), //               .startofpacket
		.output_south_endofpacket   (node_65537_output_south_endofpacket),   //               .endofpacket
		.output_south_empty         (node_65537_output_south_empty),         //               .empty
		.output_west_data           (node_65537_output_west_data),           //    output_west.data
		.output_west_valid          (node_65537_output_west_valid),          //               .valid
		.output_west_ready          (node_65537_output_west_ready),          //               .ready
		.output_west_startofpacket  (node_65537_output_west_startofpacket),  //               .startofpacket
		.output_west_endofpacket    (node_65537_output_west_endofpacket),    //               .endofpacket
		.output_west_empty          (node_65537_output_west_empty),          //               .empty
		.processing_mem_address     (node_65537_mem_address),                // processing_mem.address
		.processing_mem_readdata    (node_65537_mem_readdata),               //               .readdata
		.processing_mem_write       (node_65537_mem_write),                  //               .write
		.processing_mem_writedata   (node_65537_mem_writedata),              //               .writedata
		.reset_reset_n              (reset_reset_n)                          //          reset.reset_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_east_0 (
		.reset_n       (~rst_controller_reset_out_reset),  //  reset.reset_n
		.clk           (clk_clk),                          //  clock.clk
		.data          (node_1_output_east_data),          //     s1.data
		.empty         (node_1_output_east_empty),         //       .empty
		.endofpacket   (node_1_output_east_endofpacket),   //       .endofpacket
		.ready         (node_1_output_east_ready),         //       .ready
		.startofpacket (node_1_output_east_startofpacket), //       .startofpacket
		.valid         (node_1_output_east_valid),         //       .valid
		.readdata      (east_0_mem_readdata),              // status.readdata
		.address       (east_0_mem_address),               //       .address
		.read_n        (east_0_mem_read_n)                 //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_east_1 (
		.reset_n       (~rst_controller_reset_out_reset),      //  reset.reset_n
		.clk           (clk_clk),                              //  clock.clk
		.data          (node_65537_output_east_data),          //     s1.data
		.empty         (node_65537_output_east_empty),         //       .empty
		.endofpacket   (node_65537_output_east_endofpacket),   //       .endofpacket
		.ready         (node_65537_output_east_ready),         //       .ready
		.startofpacket (node_65537_output_east_startofpacket), //       .startofpacket
		.valid         (node_65537_output_east_valid),         //       .valid
		.readdata      (east_1_mem_readdata),                  // status.readdata
		.address       (east_1_mem_address),                   //       .address
		.read_n        (east_1_mem_read_n)                     //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_0 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_0_output_north_data),          //     s1.data
		.empty         (node_0_output_north_empty),         //       .empty
		.endofpacket   (node_0_output_north_endofpacket),   //       .endofpacket
		.ready         (node_0_output_north_ready),         //       .ready
		.startofpacket (node_0_output_north_startofpacket), //       .startofpacket
		.valid         (node_0_output_north_valid),         //       .valid
		.readdata      (north_0_mem_readdata),              // status.readdata
		.address       (north_0_mem_address),               //       .address
		.read_n        (north_0_mem_read_n)                 //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_1 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_1_output_north_data),          //     s1.data
		.empty         (node_1_output_north_empty),         //       .empty
		.endofpacket   (node_1_output_north_endofpacket),   //       .endofpacket
		.ready         (node_1_output_north_ready),         //       .ready
		.startofpacket (node_1_output_north_startofpacket), //       .startofpacket
		.valid         (node_1_output_north_valid),         //       .valid
		.readdata      (north_1_mem_readdata),              // status.readdata
		.address       (north_1_mem_address),               //       .address
		.read_n        (north_1_mem_read_n)                 //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_0 (
		.reset_n       (~rst_controller_reset_out_reset),       //  reset.reset_n
		.clk           (clk_clk),                               //  clock.clk
		.data          (node_65536_output_south_data),          //     s1.data
		.empty         (node_65536_output_south_empty),         //       .empty
		.endofpacket   (node_65536_output_south_endofpacket),   //       .endofpacket
		.ready         (node_65536_output_south_ready),         //       .ready
		.startofpacket (node_65536_output_south_startofpacket), //       .startofpacket
		.valid         (node_65536_output_south_valid),         //       .valid
		.readdata      (south_0_mem_readdata),                  // status.readdata
		.address       (south_0_mem_address),                   //       .address
		.read_n        (south_0_mem_read_n)                     //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_1 (
		.reset_n       (~rst_controller_reset_out_reset),       //  reset.reset_n
		.clk           (clk_clk),                               //  clock.clk
		.data          (node_65537_output_south_data),          //     s1.data
		.empty         (node_65537_output_south_empty),         //       .empty
		.endofpacket   (node_65537_output_south_endofpacket),   //       .endofpacket
		.ready         (node_65537_output_south_ready),         //       .ready
		.startofpacket (node_65537_output_south_startofpacket), //       .startofpacket
		.valid         (node_65537_output_south_valid),         //       .valid
		.readdata      (south_1_mem_readdata),                  // status.readdata
		.address       (south_1_mem_address),                   //       .address
		.read_n        (south_1_mem_read_n)                     //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_west_0 (
		.reset_n       (~rst_controller_reset_out_reset),  //  reset.reset_n
		.clk           (clk_clk),                          //  clock.clk
		.data          (node_0_output_west_data),          //     s1.data
		.empty         (node_0_output_west_empty),         //       .empty
		.endofpacket   (node_0_output_west_endofpacket),   //       .endofpacket
		.ready         (node_0_output_west_ready),         //       .ready
		.startofpacket (node_0_output_west_startofpacket), //       .startofpacket
		.valid         (node_0_output_west_valid),         //       .valid
		.readdata      (west_0_mem_readdata),              // status.readdata
		.address       (west_0_mem_address),               //       .address
		.read_n        (west_0_mem_read_n)                 //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_west_1 (
		.reset_n       (~rst_controller_reset_out_reset),      //  reset.reset_n
		.clk           (clk_clk),                              //  clock.clk
		.data          (node_65536_output_west_data),          //     s1.data
		.empty         (node_65536_output_west_empty),         //       .empty
		.endofpacket   (node_65536_output_west_endofpacket),   //       .endofpacket
		.ready         (node_65536_output_west_ready),         //       .ready
		.startofpacket (node_65536_output_west_startofpacket), //       .startofpacket
		.valid         (node_65536_output_west_valid),         //       .valid
		.readdata      (west_1_mem_readdata),                  // status.readdata
		.address       (west_1_mem_address),                   //       .address
		.read_n        (west_1_mem_read_n)                     //       .read_n
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
