// dircc_system_nios_single.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module dircc_system_nios_single (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         processing_stream_out_valid;         // processing:stream_out_valid -> processing:stream_in_valid
	wire  [31:0] processing_stream_out_data;          // processing:stream_out_data -> processing:stream_in_data
	wire         processing_stream_out_ready;         // processing:stream_in_ready -> processing:stream_out_ready
	wire         processing_stream_out_startofpacket; // processing:stream_out_startofpacket -> processing:stream_in_startofpacket
	wire         processing_stream_out_endofpacket;   // processing:stream_out_endofpacket -> processing:stream_in_endofpacket
	wire   [1:0] processing_stream_out_empty;         // processing:stream_out_empty -> processing:stream_in_empty
	wire  [31:0] address_address_processing_address;  // address:address_processing -> processing:address_address
	wire         rst_controller_reset_out_reset;      // rst_controller:reset_out -> [processing:reset_processing_reset_n, processing:reset_routing_reset_n]

	dircc_address_gen #(
		.ADDRESS (0)
	) address (
		.address_processing (address_address_processing_address), // address_processing.address
		.address_routing    ()                                    //    address_routing.address
	);

	dircc_system_nios_single_processing processing (
		.address_address          (address_address_processing_address),  //          address.address
		.clk_processing_clk       (clk_clk),                             //   clk_processing.clk
		.clk_routing_clk          (clk_clk),                             //      clk_routing.clk
		.mem_address              (),                                    //              mem.address
		.mem_chipselect           (),                                    //                 .chipselect
		.mem_clken                (),                                    //                 .clken
		.mem_write                (),                                    //                 .write
		.mem_readdata             (),                                    //                 .readdata
		.mem_writedata            (),                                    //                 .writedata
		.mem_byteenable           (),                                    //                 .byteenable
		.reset_processing_reset_n (~rst_controller_reset_out_reset),     // reset_processing.reset_n
		.reset_routing_reset_n    (~rst_controller_reset_out_reset),     //    reset_routing.reset_n
		.stream_in_valid          (processing_stream_out_valid),         //        stream_in.valid
		.stream_in_data           (processing_stream_out_data),          //                 .data
		.stream_in_startofpacket  (processing_stream_out_startofpacket), //                 .startofpacket
		.stream_in_endofpacket    (processing_stream_out_endofpacket),   //                 .endofpacket
		.stream_in_empty          (processing_stream_out_empty),         //                 .empty
		.stream_in_ready          (processing_stream_out_ready),         //                 .ready
		.stream_out_valid         (processing_stream_out_valid),         //       stream_out.valid
		.stream_out_data          (processing_stream_out_data),          //                 .data
		.stream_out_startofpacket (processing_stream_out_startofpacket), //                 .startofpacket
		.stream_out_endofpacket   (processing_stream_out_endofpacket),   //                 .endofpacket
		.stream_out_empty         (processing_stream_out_empty),         //                 .empty
		.stream_out_ready         (processing_stream_out_ready)          //                 .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
