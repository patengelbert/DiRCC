// dircc_status_register_tb.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_status_register_tb (
	);

	wire  [15:0] dircc_status_register_inst_mem_bfm_m0_readdata;
	wire  [15:0] dircc_status_register_inst_mem_bfm_m0_writedata;
	wire  [14:0] dircc_status_register_inst_mem_bfm_m0_address;
	wire         dircc_status_register_inst_mem_bfm_m0_write; 
	wire         dircc_status_register_inst_clk_bfm_clk_clk;          
	wire         dircc_status_register_inst_reset_bfm_reset_reset;

	dircc_status_register dircc_status_register_inst (
		.clk          	  (dircc_status_register_inst_clk_bfm_clk_clk),          //    clk.clk
		.reset_n    	  (dircc_status_register_inst_reset_bfm_reset_reset),    //  reset.reset_n
		.mem_readdata  	  (dircc_status_register_inst_mem_bfm_m0_readdata),   	 //    mem.readdata
		.mem_writedata 	  (dircc_status_register_inst_mem_bfm_m0_writedata),  	 //       .writedata
		.mem_address   	  (dircc_status_register_inst_mem_bfm_m0_address),    	 //       .address
		.mem_write     	  (dircc_status_register_inst_mem_bfm_m0_write)       	 //       .write
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dircc_status_register_inst_clk_bfm (
		.clk (dircc_status_register_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dircc_status_register_inst_reset_bfm (
		.reset (dircc_status_register_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dircc_status_register_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (15),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (2),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (0),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (0),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) dircc_status_register_inst_status_bfm (
		.clk                    (dircc_status_register_inst_clk_bfm_clk_clk),        		//       clk.clk
		.reset                  (~dircc_status_register_inst_reset_bfm_reset_reset), 		// clk_reset.reset
		.avm_address            (dircc_status_register_inst_mem_bfm_m0_address),  			//        m0.address
		.avm_readdata           (dircc_status_register_inst_mem_bfm_m0_readdata), 			//          .readdata
		.avm_writedata          (dircc_status_register_inst_mem_bfm_m0_writedata), 			//          .writedata 
		.avm_write              (dircc_status_register_inst_mem_bfm_m0_write),              // 			.write   
		.avm_read               (),     													// (terminated)
		.avm_burstcount         (),                                                         // (terminated)                             // (terminated)
		.avm_begintransfer      (),                                                         // (terminated)
		.avm_beginbursttransfer (),                                                         // (terminated)
		.avm_waitrequest        (1'b0),                                                     // (terminated)
		.avm_byteenable         (),                                                         // (terminated)
		.avm_readdatavalid      (1'b0),                                                     // (terminated)
		.avm_arbiterlock        (),                                                         // (terminated)
		.avm_lock               (),                                                         // (terminated)
		.avm_debugaccess        (),                                                         // (terminated)
		.avm_transactionid      (),                                                         // (terminated)
		.avm_readid             (8'b00000000),                                              // (terminated)
		.avm_writeid            (8'b00000000),                                              // (terminated)
		.avm_clken              (),                                                         // (terminated)
		.avm_response           (2'b00),                                                    // (terminated)
		.avm_writeresponsevalid (1'b0),                                                     // (terminated)
		.avm_writeresponserequest(),													    // (terminated)
		.avm_readresponse       (1'b0),                                                     // (terminated)
		.avm_writeresponse      (1'b0)                                                      // (terminated)
	);

endmodule
