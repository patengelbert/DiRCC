// dircc_system_node_dual.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module dircc_system_node_dual (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         node_0_output_east_valid;         // node_0:output_east_valid -> node_1:input_west_valid
	wire  [31:0] node_0_output_east_data;          // node_0:output_east_data -> node_1:input_west_data
	wire         node_0_output_east_ready;         // node_1:input_west_ready -> node_0:output_east_ready
	wire         node_0_output_east_startofpacket; // node_0:output_east_startofpacket -> node_1:input_west_startofpacket
	wire         node_0_output_east_endofpacket;   // node_0:output_east_endofpacket -> node_1:input_west_endofpacket
	wire   [1:0] node_0_output_east_empty;         // node_0:output_east_empty -> node_1:input_west_empty
	wire         node_1_output_west_valid;         // node_1:output_west_valid -> node_0:input_east_valid
	wire  [31:0] node_1_output_west_data;          // node_1:output_west_data -> node_0:input_east_data
	wire         node_1_output_west_ready;         // node_0:input_east_ready -> node_1:output_west_ready
	wire         node_1_output_west_startofpacket; // node_1:output_west_startofpacket -> node_0:input_east_startofpacket
	wire         node_1_output_west_endofpacket;   // node_1:output_west_endofpacket -> node_0:input_east_endofpacket
	wire   [1:0] node_1_output_west_empty;         // node_1:output_west_empty -> node_0:input_east_empty
	wire         rst_controller_reset_out_reset;   // rst_controller:reset_out -> [node_0:reset_processing_reset_n, node_0:reset_routing_reset_n, node_1:reset_processing_reset_n, node_1:reset_routing_reset_n]

	dircc_system_node_dual_node_0 node_0 (
		.clk_processing_clk         (clk_clk),                          //   clk_processing.clk
		.clk_routing_clk            (clk_clk),                          //      clk_routing.clk
		.input_east_data            (node_1_output_west_data),          //       input_east.data
		.input_east_valid           (node_1_output_west_valid),         //                 .valid
		.input_east_ready           (node_1_output_west_ready),         //                 .ready
		.input_east_startofpacket   (node_1_output_west_startofpacket), //                 .startofpacket
		.input_east_endofpacket     (node_1_output_west_endofpacket),   //                 .endofpacket
		.input_east_empty           (node_1_output_west_empty),         //                 .empty
		.input_north_data           (),                                 //      input_north.data
		.input_north_valid          (),                                 //                 .valid
		.input_north_ready          (),                                 //                 .ready
		.input_north_startofpacket  (),                                 //                 .startofpacket
		.input_north_endofpacket    (),                                 //                 .endofpacket
		.input_north_empty          (),                                 //                 .empty
		.input_south_data           (),                                 //      input_south.data
		.input_south_valid          (),                                 //                 .valid
		.input_south_ready          (),                                 //                 .ready
		.input_south_startofpacket  (),                                 //                 .startofpacket
		.input_south_endofpacket    (),                                 //                 .endofpacket
		.input_south_empty          (),                                 //                 .empty
		.input_west_data            (),                                 //       input_west.data
		.input_west_valid           (),                                 //                 .valid
		.input_west_ready           (),                                 //                 .ready
		.input_west_startofpacket   (),                                 //                 .startofpacket
		.input_west_endofpacket     (),                                 //                 .endofpacket
		.input_west_empty           (),                                 //                 .empty
		.output_east_data           (node_0_output_east_data),          //      output_east.data
		.output_east_valid          (node_0_output_east_valid),         //                 .valid
		.output_east_ready          (node_0_output_east_ready),         //                 .ready
		.output_east_startofpacket  (node_0_output_east_startofpacket), //                 .startofpacket
		.output_east_endofpacket    (node_0_output_east_endofpacket),   //                 .endofpacket
		.output_east_empty          (node_0_output_east_empty),         //                 .empty
		.output_north_data          (),                                 //     output_north.data
		.output_north_valid         (),                                 //                 .valid
		.output_north_ready         (),                                 //                 .ready
		.output_north_startofpacket (),                                 //                 .startofpacket
		.output_north_endofpacket   (),                                 //                 .endofpacket
		.output_north_empty         (),                                 //                 .empty
		.output_south_data          (),                                 //     output_south.data
		.output_south_valid         (),                                 //                 .valid
		.output_south_ready         (),                                 //                 .ready
		.output_south_startofpacket (),                                 //                 .startofpacket
		.output_south_endofpacket   (),                                 //                 .endofpacket
		.output_south_empty         (),                                 //                 .empty
		.output_west_data           (),                                 //      output_west.data
		.output_west_valid          (),                                 //                 .valid
		.output_west_ready          (),                                 //                 .ready
		.output_west_startofpacket  (),                                 //                 .startofpacket
		.output_west_endofpacket    (),                                 //                 .endofpacket
		.output_west_empty          (),                                 //                 .empty
		.processing_mem_address     (),                                 //   processing_mem.address
		.processing_mem_chipselect  (),                                 //                 .chipselect
		.processing_mem_clken       (),                                 //                 .clken
		.processing_mem_write       (),                                 //                 .write
		.processing_mem_readdata    (),                                 //                 .readdata
		.processing_mem_writedata   (),                                 //                 .writedata
		.processing_mem_byteenable  (),                                 //                 .byteenable
		.reset_processing_reset_n   (~rst_controller_reset_out_reset),  // reset_processing.reset_n
		.reset_routing_reset_n      (~rst_controller_reset_out_reset)   //    reset_routing.reset_n
	);

	dircc_system_node_dual_node_1 node_1 (
		.clk_processing_clk         (clk_clk),                          //   clk_processing.clk
		.clk_routing_clk            (clk_clk),                          //      clk_routing.clk
		.input_east_data            (),                                 //       input_east.data
		.input_east_valid           (),                                 //                 .valid
		.input_east_ready           (),                                 //                 .ready
		.input_east_startofpacket   (),                                 //                 .startofpacket
		.input_east_endofpacket     (),                                 //                 .endofpacket
		.input_east_empty           (),                                 //                 .empty
		.input_north_data           (),                                 //      input_north.data
		.input_north_valid          (),                                 //                 .valid
		.input_north_ready          (),                                 //                 .ready
		.input_north_startofpacket  (),                                 //                 .startofpacket
		.input_north_endofpacket    (),                                 //                 .endofpacket
		.input_north_empty          (),                                 //                 .empty
		.input_south_data           (),                                 //      input_south.data
		.input_south_valid          (),                                 //                 .valid
		.input_south_ready          (),                                 //                 .ready
		.input_south_startofpacket  (),                                 //                 .startofpacket
		.input_south_endofpacket    (),                                 //                 .endofpacket
		.input_south_empty          (),                                 //                 .empty
		.input_west_data            (node_0_output_east_data),          //       input_west.data
		.input_west_valid           (node_0_output_east_valid),         //                 .valid
		.input_west_ready           (node_0_output_east_ready),         //                 .ready
		.input_west_startofpacket   (node_0_output_east_startofpacket), //                 .startofpacket
		.input_west_endofpacket     (node_0_output_east_endofpacket),   //                 .endofpacket
		.input_west_empty           (node_0_output_east_empty),         //                 .empty
		.output_east_data           (),                                 //      output_east.data
		.output_east_valid          (),                                 //                 .valid
		.output_east_ready          (),                                 //                 .ready
		.output_east_startofpacket  (),                                 //                 .startofpacket
		.output_east_endofpacket    (),                                 //                 .endofpacket
		.output_east_empty          (),                                 //                 .empty
		.output_north_data          (),                                 //     output_north.data
		.output_north_valid         (),                                 //                 .valid
		.output_north_ready         (),                                 //                 .ready
		.output_north_startofpacket (),                                 //                 .startofpacket
		.output_north_endofpacket   (),                                 //                 .endofpacket
		.output_north_empty         (),                                 //                 .empty
		.output_south_data          (),                                 //     output_south.data
		.output_south_valid         (),                                 //                 .valid
		.output_south_ready         (),                                 //                 .ready
		.output_south_startofpacket (),                                 //                 .startofpacket
		.output_south_endofpacket   (),                                 //                 .endofpacket
		.output_south_empty         (),                                 //                 .empty
		.output_west_data           (node_1_output_west_data),          //      output_west.data
		.output_west_valid          (node_1_output_west_valid),         //                 .valid
		.output_west_ready          (node_1_output_west_ready),         //                 .ready
		.output_west_startofpacket  (node_1_output_west_startofpacket), //                 .startofpacket
		.output_west_endofpacket    (node_1_output_west_endofpacket),   //                 .endofpacket
		.output_west_empty          (node_1_output_west_empty),         //                 .empty
		.processing_mem_address     (),                                 //   processing_mem.address
		.processing_mem_chipselect  (),                                 //                 .chipselect
		.processing_mem_clken       (),                                 //                 .clken
		.processing_mem_write       (),                                 //                 .write
		.processing_mem_readdata    (),                                 //                 .readdata
		.processing_mem_writedata   (),                                 //                 .writedata
		.processing_mem_byteenable  (),                                 //                 .byteenable
		.reset_processing_reset_n   (~rst_controller_reset_out_reset),  // reset_processing.reset_n
		.reset_routing_reset_n      (~rst_controller_reset_out_reset)   //    reset_routing.reset_n
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
