// dircc_avalon_st_packet_receiver_tb.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_avalon_st_packet_receiver_tb (
	);

	import dircc_types_pkg::*;

	wire         dircc_avalon_st_packet_receiver_inst_input_valid;                 
	wire  [31:0] dircc_avalon_st_packet_receiver_inst_input_data;                  
	wire         dircc_avalon_st_packet_receiver_inst_input_ready;                 
	wire         dircc_avalon_st_packet_receiver_inst_input_startofpacket;         
	wire         dircc_avalon_st_packet_receiver_inst_input_endofpacket;           
	wire   [1:0] dircc_avalon_st_packet_receiver_inst_input_empty;
	wire         dircc_avalon_st_packet_receiver_inst_clk_bfm_clk_clk;
	wire         dircc_avalon_st_packet_receiver_inst_reset_bfm_reset_reset;
	wire         dircc_avalon_st_packet_receiver_inst_receive_done;
	wire		 dircc_avalon_st_packet_receiver_inst_receive_nearly_done;
	wire         dircc_avalon_st_packet_receiver_inst_packet_valid;
	packet_t     dircc_avalon_st_packet_receiver_inst_packet_data;
	logic 		 dircc_avalon_st_packet_receiver_inst_booting;

	dircc_avalon_st_packet_receiver dircc_avalon_st_packet_receiver_inst (
		.clk	                    (dircc_avalon_st_packet_receiver_inst_clk_bfm_clk_clk),                   //          clk.clk
		.data           			(dircc_avalon_st_packet_receiver_inst_input_data),                  	  //  	    input.data
		.valid          			(dircc_avalon_st_packet_receiver_inst_input_valid),                 	  //             .valid
		.ready          			(dircc_avalon_st_packet_receiver_inst_input_ready),                 	  //             .ready
		.startofpacket  			(dircc_avalon_st_packet_receiver_inst_input_startofpacket),         	  //             .startofpacket
		.endofpacket    			(dircc_avalon_st_packet_receiver_inst_input_endofpacket),           	  //             .endofpacket
		.empty          			(dircc_avalon_st_packet_receiver_inst_input_empty),                 	  //             .empty
		.reset_n              		(dircc_avalon_st_packet_receiver_inst_reset_bfm_reset_reset),             //        reset.reset_n
		.receive_done				(dircc_avalon_st_packet_receiver_inst_receive_done),					  //	  receive.done
		.receive_nearly_done		(dircc_avalon_st_packet_receiver_inst_receive_nearly_done),				  //             .nearly_done
		.packet_valid				(dircc_avalon_st_packet_receiver_inst_packet_valid),					  //       packet.valid
		.packet_data				(dircc_avalon_st_packet_receiver_inst_packet_data),						  //             .data
		.booting					(dircc_avalon_st_packet_receiver_inst_booting)						  	  //      booting.active
);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dircc_avalon_st_packet_receiver_inst_clk_bfm (
		.clk (dircc_avalon_st_packet_receiver_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (0),
		.VHDL_ID          (0)
	) dircc_avalon_st_packet_receiver_inst_input_bfm (
		.clk                (dircc_avalon_st_packet_receiver_inst_clk_bfm_clk_clk),         //       clk.clk
		.reset              (~dircc_avalon_st_packet_receiver_inst_reset_bfm_reset_reset),  // clk_reset.reset
		.src_data           (dircc_avalon_st_packet_receiver_inst_input_data),          	//       src.data
		.src_valid          (dircc_avalon_st_packet_receiver_inst_input_valid),         	//          .valid
		.src_ready          (dircc_avalon_st_packet_receiver_inst_input_ready),         	//          .ready
		.src_startofpacket  (dircc_avalon_st_packet_receiver_inst_input_startofpacket), 	//          .startofpacket
		.src_endofpacket    (dircc_avalon_st_packet_receiver_inst_input_endofpacket),   	//          .endofpacket
		.src_empty          (dircc_avalon_st_packet_receiver_inst_input_empty),         	//          .empty
		.src_channel        (),                                         					// (terminated)
		.src_error          ()                                          					// (terminated)
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dircc_avalon_st_packet_receiver_inst_reset_bfm (
		.reset (dircc_avalon_st_packet_receiver_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dircc_avalon_st_packet_receiver_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
