// test.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module test (
		input  wire        clk_clk,                                   //                         clk.clk
		input  wire        reset_reset_n,                             //                       reset.reset_n
		output wire        st_pipeline_stage_0_sink0_ready,           //   st_pipeline_stage_0_sink0.ready
		input  wire        st_pipeline_stage_0_sink0_valid,           //                            .valid
		input  wire        st_pipeline_stage_0_sink0_startofpacket,   //                            .startofpacket
		input  wire        st_pipeline_stage_0_sink0_endofpacket,     //                            .endofpacket
		input  wire [31:0] st_pipeline_stage_0_sink0_data,            //                            .data
		input  wire        st_pipeline_stage_0_source0_ready,         // st_pipeline_stage_0_source0.ready
		output wire        st_pipeline_stage_0_source0_valid,         //                            .valid
		output wire        st_pipeline_stage_0_source0_startofpacket, //                            .startofpacket
		output wire        st_pipeline_stage_0_source0_endofpacket,   //                            .endofpacket
		output wire [31:0] st_pipeline_stage_0_source0_data           //                            .data
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> st_pipeline_stage_0:reset

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (4),
		.BITS_PER_SYMBOL  (8),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) st_pipeline_stage_0 (
		.clk               (clk_clk),                                   //       cr0.clk
		.reset             (rst_controller_reset_out_reset),            // cr0_reset.reset
		.in_ready          (st_pipeline_stage_0_sink0_ready),           //     sink0.ready
		.in_valid          (st_pipeline_stage_0_sink0_valid),           //          .valid
		.in_startofpacket  (st_pipeline_stage_0_sink0_startofpacket),   //          .startofpacket
		.in_endofpacket    (st_pipeline_stage_0_sink0_endofpacket),     //          .endofpacket
		.in_data           (st_pipeline_stage_0_sink0_data),            //          .data
		.out_ready         (st_pipeline_stage_0_source0_ready),         //   source0.ready
		.out_valid         (st_pipeline_stage_0_source0_valid),         //          .valid
		.out_startofpacket (st_pipeline_stage_0_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (st_pipeline_stage_0_source0_endofpacket),   //          .endofpacket
		.out_data          (st_pipeline_stage_0_source0_data),          //          .data
		.in_empty          (1'b0),                                      // (terminated)
		.out_empty         (),                                          // (terminated)
		.out_error         (),                                          // (terminated)
		.in_error          (1'b0),                                      // (terminated)
		.out_channel       (),                                          // (terminated)
		.in_channel        (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
