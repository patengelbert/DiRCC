// demo.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module demo (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         streaming_0_stream_out_valid;         // streaming_0:stream_out_valid -> streaming_0:stream_in_valid
	wire  [31:0] streaming_0_stream_out_data;          // streaming_0:stream_out_data -> streaming_0:stream_in_data
	wire         streaming_0_stream_out_ready;         // streaming_0:stream_in_ready -> streaming_0:stream_out_ready
	wire         streaming_0_stream_out_startofpacket; // streaming_0:stream_out_startofpacket -> streaming_0:stream_in_startofpacket
	wire         streaming_0_stream_out_endofpacket;   // streaming_0:stream_out_endofpacket -> streaming_0:stream_in_endofpacket
	wire   [1:0] streaming_0_stream_out_empty;         // streaming_0:stream_out_empty -> streaming_0:stream_in_empty

	demo_streaming_0 streaming_0 (
		.clk_clk                  (clk_clk),                              //        clk.clk
		.reset_reset_n            (reset_reset_n),                        //      reset.reset_n
		.stream_in_valid          (streaming_0_stream_out_valid),         //  stream_in.valid
		.stream_in_data           (streaming_0_stream_out_data),          //           .data
		.stream_in_startofpacket  (streaming_0_stream_out_startofpacket), //           .startofpacket
		.stream_in_endofpacket    (streaming_0_stream_out_endofpacket),   //           .endofpacket
		.stream_in_empty          (streaming_0_stream_out_empty),         //           .empty
		.stream_in_ready          (streaming_0_stream_out_ready),         //           .ready
		.stream_out_valid         (streaming_0_stream_out_valid),         // stream_out.valid
		.stream_out_data          (streaming_0_stream_out_data),          //           .data
		.stream_out_startofpacket (streaming_0_stream_out_startofpacket), //           .startofpacket
		.stream_out_endofpacket   (streaming_0_stream_out_endofpacket),   //           .endofpacket
		.stream_out_empty         (streaming_0_stream_out_empty),         //           .empty
		.stream_out_ready         (streaming_0_stream_out_ready)          //           .ready
	);

endmodule
