// dircc_system_nios_single.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module dircc_system_nios_single (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         node_0_stream_out_valid;         // node_0:stream_out_valid -> node_0:stream_in_valid
	wire  [31:0] node_0_stream_out_data;          // node_0:stream_out_data -> node_0:stream_in_data
	wire         node_0_stream_out_ready;         // node_0:stream_in_ready -> node_0:stream_out_ready
	wire         node_0_stream_out_startofpacket; // node_0:stream_out_startofpacket -> node_0:stream_in_startofpacket
	wire         node_0_stream_out_endofpacket;   // node_0:stream_out_endofpacket -> node_0:stream_in_endofpacket
	wire   [1:0] node_0_stream_out_empty;         // node_0:stream_out_empty -> node_0:stream_in_empty

	dircc_system_nios_single_node_0 node_0 (
		.clk_clk                  (clk_clk),                         //        clk.clk
		.reset_reset_n            (reset_reset_n),                   //      reset.reset_n
		.stream_in_valid          (node_0_stream_out_valid),         //  stream_in.valid
		.stream_in_data           (node_0_stream_out_data),          //           .data
		.stream_in_startofpacket  (node_0_stream_out_startofpacket), //           .startofpacket
		.stream_in_endofpacket    (node_0_stream_out_endofpacket),   //           .endofpacket
		.stream_in_empty          (node_0_stream_out_empty),         //           .empty
		.stream_in_ready          (node_0_stream_out_ready),         //           .ready
		.stream_out_valid         (node_0_stream_out_valid),         // stream_out.valid
		.stream_out_data          (node_0_stream_out_data),          //           .data
		.stream_out_startofpacket (node_0_stream_out_startofpacket), //           .startofpacket
		.stream_out_endofpacket   (node_0_stream_out_endofpacket),   //           .endofpacket
		.stream_out_empty         (node_0_stream_out_empty),         //           .empty
		.stream_out_ready         (node_0_stream_out_ready)          //           .ready
	);

endmodule
