// dircc_system_node_dual_hps.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_system_node_dual_hps (
		input  wire        clk_clk,                        //    clk.clk
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53, // hps_io.hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54, //       .hps_io_gpio_inst_GPIO54
		output wire [14:0] memory_mem_a,                   // memory.mem_a
		output wire [2:0]  memory_mem_ba,                  //       .mem_ba
		output wire        memory_mem_ck,                  //       .mem_ck
		output wire        memory_mem_ck_n,                //       .mem_ck_n
		output wire        memory_mem_cke,                 //       .mem_cke
		output wire        memory_mem_cs_n,                //       .mem_cs_n
		output wire        memory_mem_ras_n,               //       .mem_ras_n
		output wire        memory_mem_cas_n,               //       .mem_cas_n
		output wire        memory_mem_we_n,                //       .mem_we_n
		output wire        memory_mem_reset_n,             //       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                  //       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                 //       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,               //       .mem_dqs_n
		output wire        memory_mem_odt,                 //       .mem_odt
		output wire [3:0]  memory_mem_dm,                  //       .mem_dm
		input  wire        memory_oct_rzqin,               //       .oct_rzqin
		input  wire        reset_reset_n                   //  reset.reset_n
	);

	wire         node_0_output_east_valid;                           // node_0:output_east_valid -> node_1:input_west_valid
	wire  [31:0] node_0_output_east_data;                            // node_0:output_east_data -> node_1:input_west_data
	wire         node_0_output_east_ready;                           // node_1:input_west_ready -> node_0:output_east_ready
	wire         node_0_output_east_startofpacket;                   // node_0:output_east_startofpacket -> node_1:input_west_startofpacket
	wire         node_0_output_east_endofpacket;                     // node_0:output_east_endofpacket -> node_1:input_west_endofpacket
	wire   [1:0] node_0_output_east_empty;                           // node_0:output_east_empty -> node_1:input_west_empty
	wire         node_1_output_west_valid;                           // node_1:output_west_valid -> node_0:input_east_valid
	wire  [31:0] node_1_output_west_data;                            // node_1:output_west_data -> node_0:input_east_data
	wire         node_1_output_west_ready;                           // node_0:input_east_ready -> node_1:output_west_ready
	wire         node_1_output_west_startofpacket;                   // node_1:output_west_startofpacket -> node_0:input_east_startofpacket
	wire         node_1_output_west_endofpacket;                     // node_1:output_west_endofpacket -> node_0:input_east_endofpacket
	wire   [1:0] node_1_output_west_empty;                           // node_1:output_west_empty -> node_0:input_east_empty
	wire   [1:0] hps_h2f_axi_master_awburst;                         // HPS:h2f_AWBURST -> mm_interconnect_0:HPS_h2f_axi_master_awburst
	wire   [3:0] hps_h2f_axi_master_arlen;                           // HPS:h2f_ARLEN -> mm_interconnect_0:HPS_h2f_axi_master_arlen
	wire   [3:0] hps_h2f_axi_master_wstrb;                           // HPS:h2f_WSTRB -> mm_interconnect_0:HPS_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_wready;                          // mm_interconnect_0:HPS_h2f_axi_master_wready -> HPS:h2f_WREADY
	wire  [11:0] hps_h2f_axi_master_rid;                             // mm_interconnect_0:HPS_h2f_axi_master_rid -> HPS:h2f_RID
	wire         hps_h2f_axi_master_rready;                          // HPS:h2f_RREADY -> mm_interconnect_0:HPS_h2f_axi_master_rready
	wire   [3:0] hps_h2f_axi_master_awlen;                           // HPS:h2f_AWLEN -> mm_interconnect_0:HPS_h2f_axi_master_awlen
	wire  [11:0] hps_h2f_axi_master_wid;                             // HPS:h2f_WID -> mm_interconnect_0:HPS_h2f_axi_master_wid
	wire   [3:0] hps_h2f_axi_master_arcache;                         // HPS:h2f_ARCACHE -> mm_interconnect_0:HPS_h2f_axi_master_arcache
	wire         hps_h2f_axi_master_wvalid;                          // HPS:h2f_WVALID -> mm_interconnect_0:HPS_h2f_axi_master_wvalid
	wire  [29:0] hps_h2f_axi_master_araddr;                          // HPS:h2f_ARADDR -> mm_interconnect_0:HPS_h2f_axi_master_araddr
	wire   [2:0] hps_h2f_axi_master_arprot;                          // HPS:h2f_ARPROT -> mm_interconnect_0:HPS_h2f_axi_master_arprot
	wire   [2:0] hps_h2f_axi_master_awprot;                          // HPS:h2f_AWPROT -> mm_interconnect_0:HPS_h2f_axi_master_awprot
	wire  [31:0] hps_h2f_axi_master_wdata;                           // HPS:h2f_WDATA -> mm_interconnect_0:HPS_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_arvalid;                         // HPS:h2f_ARVALID -> mm_interconnect_0:HPS_h2f_axi_master_arvalid
	wire   [3:0] hps_h2f_axi_master_awcache;                         // HPS:h2f_AWCACHE -> mm_interconnect_0:HPS_h2f_axi_master_awcache
	wire  [11:0] hps_h2f_axi_master_arid;                            // HPS:h2f_ARID -> mm_interconnect_0:HPS_h2f_axi_master_arid
	wire   [1:0] hps_h2f_axi_master_arlock;                          // HPS:h2f_ARLOCK -> mm_interconnect_0:HPS_h2f_axi_master_arlock
	wire   [1:0] hps_h2f_axi_master_awlock;                          // HPS:h2f_AWLOCK -> mm_interconnect_0:HPS_h2f_axi_master_awlock
	wire  [29:0] hps_h2f_axi_master_awaddr;                          // HPS:h2f_AWADDR -> mm_interconnect_0:HPS_h2f_axi_master_awaddr
	wire   [1:0] hps_h2f_axi_master_bresp;                           // mm_interconnect_0:HPS_h2f_axi_master_bresp -> HPS:h2f_BRESP
	wire         hps_h2f_axi_master_arready;                         // mm_interconnect_0:HPS_h2f_axi_master_arready -> HPS:h2f_ARREADY
	wire  [31:0] hps_h2f_axi_master_rdata;                           // mm_interconnect_0:HPS_h2f_axi_master_rdata -> HPS:h2f_RDATA
	wire         hps_h2f_axi_master_awready;                         // mm_interconnect_0:HPS_h2f_axi_master_awready -> HPS:h2f_AWREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                         // HPS:h2f_ARBURST -> mm_interconnect_0:HPS_h2f_axi_master_arburst
	wire   [2:0] hps_h2f_axi_master_arsize;                          // HPS:h2f_ARSIZE -> mm_interconnect_0:HPS_h2f_axi_master_arsize
	wire         hps_h2f_axi_master_bready;                          // HPS:h2f_BREADY -> mm_interconnect_0:HPS_h2f_axi_master_bready
	wire         hps_h2f_axi_master_rlast;                           // mm_interconnect_0:HPS_h2f_axi_master_rlast -> HPS:h2f_RLAST
	wire         hps_h2f_axi_master_wlast;                           // HPS:h2f_WLAST -> mm_interconnect_0:HPS_h2f_axi_master_wlast
	wire   [1:0] hps_h2f_axi_master_rresp;                           // mm_interconnect_0:HPS_h2f_axi_master_rresp -> HPS:h2f_RRESP
	wire  [11:0] hps_h2f_axi_master_awid;                            // HPS:h2f_AWID -> mm_interconnect_0:HPS_h2f_axi_master_awid
	wire  [11:0] hps_h2f_axi_master_bid;                             // mm_interconnect_0:HPS_h2f_axi_master_bid -> HPS:h2f_BID
	wire         hps_h2f_axi_master_bvalid;                          // mm_interconnect_0:HPS_h2f_axi_master_bvalid -> HPS:h2f_BVALID
	wire   [2:0] hps_h2f_axi_master_awsize;                          // HPS:h2f_AWSIZE -> mm_interconnect_0:HPS_h2f_axi_master_awsize
	wire         hps_h2f_axi_master_awvalid;                         // HPS:h2f_AWVALID -> mm_interconnect_0:HPS_h2f_axi_master_awvalid
	wire         hps_h2f_axi_master_rvalid;                          // mm_interconnect_0:HPS_h2f_axi_master_rvalid -> HPS:h2f_RVALID
	wire         mm_interconnect_0_node_0_processing_mem_chipselect; // mm_interconnect_0:node_0_processing_mem_chipselect -> node_0:processing_mem_chipselect
	wire  [15:0] mm_interconnect_0_node_0_processing_mem_readdata;   // node_0:processing_mem_readdata -> mm_interconnect_0:node_0_processing_mem_readdata
	wire  [14:0] mm_interconnect_0_node_0_processing_mem_address;    // mm_interconnect_0:node_0_processing_mem_address -> node_0:processing_mem_address
	wire   [1:0] mm_interconnect_0_node_0_processing_mem_byteenable; // mm_interconnect_0:node_0_processing_mem_byteenable -> node_0:processing_mem_byteenable
	wire         mm_interconnect_0_node_0_processing_mem_write;      // mm_interconnect_0:node_0_processing_mem_write -> node_0:processing_mem_write
	wire  [15:0] mm_interconnect_0_node_0_processing_mem_writedata;  // mm_interconnect_0:node_0_processing_mem_writedata -> node_0:processing_mem_writedata
	wire         mm_interconnect_0_node_0_processing_mem_clken;      // mm_interconnect_0:node_0_processing_mem_clken -> node_0:processing_mem_clken
	wire         mm_interconnect_0_node_1_processing_mem_chipselect; // mm_interconnect_0:node_1_processing_mem_chipselect -> node_1:processing_mem_chipselect
	wire  [15:0] mm_interconnect_0_node_1_processing_mem_readdata;   // node_1:processing_mem_readdata -> mm_interconnect_0:node_1_processing_mem_readdata
	wire  [14:0] mm_interconnect_0_node_1_processing_mem_address;    // mm_interconnect_0:node_1_processing_mem_address -> node_1:processing_mem_address
	wire   [1:0] mm_interconnect_0_node_1_processing_mem_byteenable; // mm_interconnect_0:node_1_processing_mem_byteenable -> node_1:processing_mem_byteenable
	wire         mm_interconnect_0_node_1_processing_mem_write;      // mm_interconnect_0:node_1_processing_mem_write -> node_1:processing_mem_write
	wire  [15:0] mm_interconnect_0_node_1_processing_mem_writedata;  // mm_interconnect_0:node_1_processing_mem_writedata -> node_1:processing_mem_writedata
	wire         mm_interconnect_0_node_1_processing_mem_clken;      // mm_interconnect_0:node_1_processing_mem_clken -> node_1:processing_mem_clken
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [mm_interconnect_0:node_0_reset_processing_reset_bridge_in_reset_reset, node_0:reset_processing_reset_n, node_0:reset_routing_reset_n, node_1:reset_processing_reset_n, node_1:reset_routing_reset_n]
	wire         hps_h2f_reset_reset;                                // HPS:h2f_rst_n -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> mm_interconnect_0:HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	dircc_system_node_dual_hps_HPS #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps (
		.mem_a                   (memory_mem_a),                   //         memory.mem_a
		.mem_ba                  (memory_mem_ba),                  //               .mem_ba
		.mem_ck                  (memory_mem_ck),                  //               .mem_ck
		.mem_ck_n                (memory_mem_ck_n),                //               .mem_ck_n
		.mem_cke                 (memory_mem_cke),                 //               .mem_cke
		.mem_cs_n                (memory_mem_cs_n),                //               .mem_cs_n
		.mem_ras_n               (memory_mem_ras_n),               //               .mem_ras_n
		.mem_cas_n               (memory_mem_cas_n),               //               .mem_cas_n
		.mem_we_n                (memory_mem_we_n),                //               .mem_we_n
		.mem_reset_n             (memory_mem_reset_n),             //               .mem_reset_n
		.mem_dq                  (memory_mem_dq),                  //               .mem_dq
		.mem_dqs                 (memory_mem_dqs),                 //               .mem_dqs
		.mem_dqs_n               (memory_mem_dqs_n),               //               .mem_dqs_n
		.mem_odt                 (memory_mem_odt),                 //               .mem_odt
		.mem_dm                  (memory_mem_dm),                  //               .mem_dm
		.oct_rzqin               (memory_oct_rzqin),               //               .oct_rzqin
		.hps_io_gpio_inst_GPIO53 (hps_io_hps_io_gpio_inst_GPIO53), //         hps_io.hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54 (hps_io_hps_io_gpio_inst_GPIO54), //               .hps_io_gpio_inst_GPIO54
		.h2f_rst_n               (hps_h2f_reset_reset),            //      h2f_reset.reset_n
		.h2f_axi_clk             (clk_clk),                        //  h2f_axi_clock.clk
		.h2f_AWID                (hps_h2f_axi_master_awid),        // h2f_axi_master.awid
		.h2f_AWADDR              (hps_h2f_axi_master_awaddr),      //               .awaddr
		.h2f_AWLEN               (hps_h2f_axi_master_awlen),       //               .awlen
		.h2f_AWSIZE              (hps_h2f_axi_master_awsize),      //               .awsize
		.h2f_AWBURST             (hps_h2f_axi_master_awburst),     //               .awburst
		.h2f_AWLOCK              (hps_h2f_axi_master_awlock),      //               .awlock
		.h2f_AWCACHE             (hps_h2f_axi_master_awcache),     //               .awcache
		.h2f_AWPROT              (hps_h2f_axi_master_awprot),      //               .awprot
		.h2f_AWVALID             (hps_h2f_axi_master_awvalid),     //               .awvalid
		.h2f_AWREADY             (hps_h2f_axi_master_awready),     //               .awready
		.h2f_WID                 (hps_h2f_axi_master_wid),         //               .wid
		.h2f_WDATA               (hps_h2f_axi_master_wdata),       //               .wdata
		.h2f_WSTRB               (hps_h2f_axi_master_wstrb),       //               .wstrb
		.h2f_WLAST               (hps_h2f_axi_master_wlast),       //               .wlast
		.h2f_WVALID              (hps_h2f_axi_master_wvalid),      //               .wvalid
		.h2f_WREADY              (hps_h2f_axi_master_wready),      //               .wready
		.h2f_BID                 (hps_h2f_axi_master_bid),         //               .bid
		.h2f_BRESP               (hps_h2f_axi_master_bresp),       //               .bresp
		.h2f_BVALID              (hps_h2f_axi_master_bvalid),      //               .bvalid
		.h2f_BREADY              (hps_h2f_axi_master_bready),      //               .bready
		.h2f_ARID                (hps_h2f_axi_master_arid),        //               .arid
		.h2f_ARADDR              (hps_h2f_axi_master_araddr),      //               .araddr
		.h2f_ARLEN               (hps_h2f_axi_master_arlen),       //               .arlen
		.h2f_ARSIZE              (hps_h2f_axi_master_arsize),      //               .arsize
		.h2f_ARBURST             (hps_h2f_axi_master_arburst),     //               .arburst
		.h2f_ARLOCK              (hps_h2f_axi_master_arlock),      //               .arlock
		.h2f_ARCACHE             (hps_h2f_axi_master_arcache),     //               .arcache
		.h2f_ARPROT              (hps_h2f_axi_master_arprot),      //               .arprot
		.h2f_ARVALID             (hps_h2f_axi_master_arvalid),     //               .arvalid
		.h2f_ARREADY             (hps_h2f_axi_master_arready),     //               .arready
		.h2f_RID                 (hps_h2f_axi_master_rid),         //               .rid
		.h2f_RDATA               (hps_h2f_axi_master_rdata),       //               .rdata
		.h2f_RRESP               (hps_h2f_axi_master_rresp),       //               .rresp
		.h2f_RLAST               (hps_h2f_axi_master_rlast),       //               .rlast
		.h2f_RVALID              (hps_h2f_axi_master_rvalid),      //               .rvalid
		.h2f_RREADY              (hps_h2f_axi_master_rready)       //               .rready
	);

	dircc_system_node_dual_hps_node_0 node_0 (
		.clk_processing_clk         (clk_clk),                                            //   clk_processing.clk
		.clk_routing_clk            (clk_clk),                                            //      clk_routing.clk
		.input_east_data            (node_1_output_west_data),                            //       input_east.data
		.input_east_valid           (node_1_output_west_valid),                           //                 .valid
		.input_east_ready           (node_1_output_west_ready),                           //                 .ready
		.input_east_startofpacket   (node_1_output_west_startofpacket),                   //                 .startofpacket
		.input_east_endofpacket     (node_1_output_west_endofpacket),                     //                 .endofpacket
		.input_east_empty           (node_1_output_west_empty),                           //                 .empty
		.input_north_data           (),                                                   //      input_north.data
		.input_north_valid          (),                                                   //                 .valid
		.input_north_ready          (),                                                   //                 .ready
		.input_north_startofpacket  (),                                                   //                 .startofpacket
		.input_north_endofpacket    (),                                                   //                 .endofpacket
		.input_north_empty          (),                                                   //                 .empty
		.input_south_data           (),                                                   //      input_south.data
		.input_south_valid          (),                                                   //                 .valid
		.input_south_ready          (),                                                   //                 .ready
		.input_south_startofpacket  (),                                                   //                 .startofpacket
		.input_south_endofpacket    (),                                                   //                 .endofpacket
		.input_south_empty          (),                                                   //                 .empty
		.input_west_data            (),                                                   //       input_west.data
		.input_west_valid           (),                                                   //                 .valid
		.input_west_ready           (),                                                   //                 .ready
		.input_west_startofpacket   (),                                                   //                 .startofpacket
		.input_west_endofpacket     (),                                                   //                 .endofpacket
		.input_west_empty           (),                                                   //                 .empty
		.output_east_data           (node_0_output_east_data),                            //      output_east.data
		.output_east_valid          (node_0_output_east_valid),                           //                 .valid
		.output_east_ready          (node_0_output_east_ready),                           //                 .ready
		.output_east_startofpacket  (node_0_output_east_startofpacket),                   //                 .startofpacket
		.output_east_endofpacket    (node_0_output_east_endofpacket),                     //                 .endofpacket
		.output_east_empty          (node_0_output_east_empty),                           //                 .empty
		.output_north_data          (),                                                   //     output_north.data
		.output_north_valid         (),                                                   //                 .valid
		.output_north_ready         (),                                                   //                 .ready
		.output_north_startofpacket (),                                                   //                 .startofpacket
		.output_north_endofpacket   (),                                                   //                 .endofpacket
		.output_north_empty         (),                                                   //                 .empty
		.output_south_data          (),                                                   //     output_south.data
		.output_south_valid         (),                                                   //                 .valid
		.output_south_ready         (),                                                   //                 .ready
		.output_south_startofpacket (),                                                   //                 .startofpacket
		.output_south_endofpacket   (),                                                   //                 .endofpacket
		.output_south_empty         (),                                                   //                 .empty
		.output_west_data           (),                                                   //      output_west.data
		.output_west_valid          (),                                                   //                 .valid
		.output_west_ready          (),                                                   //                 .ready
		.output_west_startofpacket  (),                                                   //                 .startofpacket
		.output_west_endofpacket    (),                                                   //                 .endofpacket
		.output_west_empty          (),                                                   //                 .empty
		.processing_mem_address     (mm_interconnect_0_node_0_processing_mem_address),    //   processing_mem.address
		.processing_mem_chipselect  (mm_interconnect_0_node_0_processing_mem_chipselect), //                 .chipselect
		.processing_mem_clken       (mm_interconnect_0_node_0_processing_mem_clken),      //                 .clken
		.processing_mem_write       (mm_interconnect_0_node_0_processing_mem_write),      //                 .write
		.processing_mem_readdata    (mm_interconnect_0_node_0_processing_mem_readdata),   //                 .readdata
		.processing_mem_writedata   (mm_interconnect_0_node_0_processing_mem_writedata),  //                 .writedata
		.processing_mem_byteenable  (mm_interconnect_0_node_0_processing_mem_byteenable), //                 .byteenable
		.reset_processing_reset_n   (~rst_controller_reset_out_reset),                    // reset_processing.reset_n
		.reset_routing_reset_n      (~rst_controller_reset_out_reset)                     //    reset_routing.reset_n
	);

	dircc_system_node_dual_hps_node_1 node_1 (
		.clk_processing_clk         (clk_clk),                                            //   clk_processing.clk
		.clk_routing_clk            (clk_clk),                                            //      clk_routing.clk
		.input_east_data            (),                                                   //       input_east.data
		.input_east_valid           (),                                                   //                 .valid
		.input_east_ready           (),                                                   //                 .ready
		.input_east_startofpacket   (),                                                   //                 .startofpacket
		.input_east_endofpacket     (),                                                   //                 .endofpacket
		.input_east_empty           (),                                                   //                 .empty
		.input_north_data           (),                                                   //      input_north.data
		.input_north_valid          (),                                                   //                 .valid
		.input_north_ready          (),                                                   //                 .ready
		.input_north_startofpacket  (),                                                   //                 .startofpacket
		.input_north_endofpacket    (),                                                   //                 .endofpacket
		.input_north_empty          (),                                                   //                 .empty
		.input_south_data           (),                                                   //      input_south.data
		.input_south_valid          (),                                                   //                 .valid
		.input_south_ready          (),                                                   //                 .ready
		.input_south_startofpacket  (),                                                   //                 .startofpacket
		.input_south_endofpacket    (),                                                   //                 .endofpacket
		.input_south_empty          (),                                                   //                 .empty
		.input_west_data            (node_0_output_east_data),                            //       input_west.data
		.input_west_valid           (node_0_output_east_valid),                           //                 .valid
		.input_west_ready           (node_0_output_east_ready),                           //                 .ready
		.input_west_startofpacket   (node_0_output_east_startofpacket),                   //                 .startofpacket
		.input_west_endofpacket     (node_0_output_east_endofpacket),                     //                 .endofpacket
		.input_west_empty           (node_0_output_east_empty),                           //                 .empty
		.output_east_data           (),                                                   //      output_east.data
		.output_east_valid          (),                                                   //                 .valid
		.output_east_ready          (),                                                   //                 .ready
		.output_east_startofpacket  (),                                                   //                 .startofpacket
		.output_east_endofpacket    (),                                                   //                 .endofpacket
		.output_east_empty          (),                                                   //                 .empty
		.output_north_data          (),                                                   //     output_north.data
		.output_north_valid         (),                                                   //                 .valid
		.output_north_ready         (),                                                   //                 .ready
		.output_north_startofpacket (),                                                   //                 .startofpacket
		.output_north_endofpacket   (),                                                   //                 .endofpacket
		.output_north_empty         (),                                                   //                 .empty
		.output_south_data          (),                                                   //     output_south.data
		.output_south_valid         (),                                                   //                 .valid
		.output_south_ready         (),                                                   //                 .ready
		.output_south_startofpacket (),                                                   //                 .startofpacket
		.output_south_endofpacket   (),                                                   //                 .endofpacket
		.output_south_empty         (),                                                   //                 .empty
		.output_west_data           (node_1_output_west_data),                            //      output_west.data
		.output_west_valid          (node_1_output_west_valid),                           //                 .valid
		.output_west_ready          (node_1_output_west_ready),                           //                 .ready
		.output_west_startofpacket  (node_1_output_west_startofpacket),                   //                 .startofpacket
		.output_west_endofpacket    (node_1_output_west_endofpacket),                     //                 .endofpacket
		.output_west_empty          (node_1_output_west_empty),                           //                 .empty
		.processing_mem_address     (mm_interconnect_0_node_1_processing_mem_address),    //   processing_mem.address
		.processing_mem_chipselect  (mm_interconnect_0_node_1_processing_mem_chipselect), //                 .chipselect
		.processing_mem_clken       (mm_interconnect_0_node_1_processing_mem_clken),      //                 .clken
		.processing_mem_write       (mm_interconnect_0_node_1_processing_mem_write),      //                 .write
		.processing_mem_readdata    (mm_interconnect_0_node_1_processing_mem_readdata),   //                 .readdata
		.processing_mem_writedata   (mm_interconnect_0_node_1_processing_mem_writedata),  //                 .writedata
		.processing_mem_byteenable  (mm_interconnect_0_node_1_processing_mem_byteenable), //                 .byteenable
		.reset_processing_reset_n   (~rst_controller_reset_out_reset),                    // reset_processing.reset_n
		.reset_routing_reset_n      (~rst_controller_reset_out_reset)                     //    reset_routing.reset_n
	);

	dircc_system_node_dual_hps_mm_interconnect_0 mm_interconnect_0 (
		.HPS_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),                            //                                       HPS_h2f_axi_master.awid
		.HPS_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),                          //                                                         .awaddr
		.HPS_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),                           //                                                         .awlen
		.HPS_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),                          //                                                         .awsize
		.HPS_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),                         //                                                         .awburst
		.HPS_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),                          //                                                         .awlock
		.HPS_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),                         //                                                         .awcache
		.HPS_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),                          //                                                         .awprot
		.HPS_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),                         //                                                         .awvalid
		.HPS_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),                         //                                                         .awready
		.HPS_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),                             //                                                         .wid
		.HPS_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),                           //                                                         .wdata
		.HPS_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),                           //                                                         .wstrb
		.HPS_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),                           //                                                         .wlast
		.HPS_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),                          //                                                         .wvalid
		.HPS_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),                          //                                                         .wready
		.HPS_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),                             //                                                         .bid
		.HPS_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),                           //                                                         .bresp
		.HPS_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),                          //                                                         .bvalid
		.HPS_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),                          //                                                         .bready
		.HPS_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),                            //                                                         .arid
		.HPS_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),                          //                                                         .araddr
		.HPS_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),                           //                                                         .arlen
		.HPS_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),                          //                                                         .arsize
		.HPS_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),                         //                                                         .arburst
		.HPS_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),                          //                                                         .arlock
		.HPS_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),                         //                                                         .arcache
		.HPS_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),                          //                                                         .arprot
		.HPS_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),                         //                                                         .arvalid
		.HPS_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),                         //                                                         .arready
		.HPS_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),                             //                                                         .rid
		.HPS_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),                           //                                                         .rdata
		.HPS_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),                           //                                                         .rresp
		.HPS_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),                           //                                                         .rlast
		.HPS_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),                          //                                                         .rvalid
		.HPS_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),                          //                                                         .rready
		.clk_clk_clk                                                    (clk_clk),                                            //                                                  clk_clk.clk
		.HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                 // HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.node_0_reset_processing_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                     //            node_0_reset_processing_reset_bridge_in_reset.reset
		.node_0_processing_mem_address                                  (mm_interconnect_0_node_0_processing_mem_address),    //                                    node_0_processing_mem.address
		.node_0_processing_mem_write                                    (mm_interconnect_0_node_0_processing_mem_write),      //                                                         .write
		.node_0_processing_mem_readdata                                 (mm_interconnect_0_node_0_processing_mem_readdata),   //                                                         .readdata
		.node_0_processing_mem_writedata                                (mm_interconnect_0_node_0_processing_mem_writedata),  //                                                         .writedata
		.node_0_processing_mem_byteenable                               (mm_interconnect_0_node_0_processing_mem_byteenable), //                                                         .byteenable
		.node_0_processing_mem_chipselect                               (mm_interconnect_0_node_0_processing_mem_chipselect), //                                                         .chipselect
		.node_0_processing_mem_clken                                    (mm_interconnect_0_node_0_processing_mem_clken),      //                                                         .clken
		.node_1_processing_mem_address                                  (mm_interconnect_0_node_1_processing_mem_address),    //                                    node_1_processing_mem.address
		.node_1_processing_mem_write                                    (mm_interconnect_0_node_1_processing_mem_write),      //                                                         .write
		.node_1_processing_mem_readdata                                 (mm_interconnect_0_node_1_processing_mem_readdata),   //                                                         .readdata
		.node_1_processing_mem_writedata                                (mm_interconnect_0_node_1_processing_mem_writedata),  //                                                         .writedata
		.node_1_processing_mem_byteenable                               (mm_interconnect_0_node_1_processing_mem_byteenable), //                                                         .byteenable
		.node_1_processing_mem_chipselect                               (mm_interconnect_0_node_1_processing_mem_chipselect), //                                                         .chipselect
		.node_1_processing_mem_clken                                    (mm_interconnect_0_node_1_processing_mem_clken)       //                                                         .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (~hps_h2f_reset_reset),           // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
