// dircc_system_rtl_gals_test_version.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module dircc_system_rtl_gals_test_version (
		input  wire        clk_clk,                   //             clk.clk
		input  wire [14:0] node_0_mem_address,        //      node_0_mem.address
		output wire [15:0] node_0_mem_readdata,       //                .readdata
		input  wire        node_0_mem_write,          //                .write
		input  wire [15:0] node_0_mem_writedata,      //                .writedata
		input  wire [14:0] node_131072_mem_address,   // node_131072_mem.address
		output wire [15:0] node_131072_mem_readdata,  //                .readdata
		input  wire        node_131072_mem_write,     //                .write
		input  wire [15:0] node_131072_mem_writedata, //                .writedata
		input  wire [14:0] node_131073_mem_address,   // node_131073_mem.address
		output wire [15:0] node_131073_mem_readdata,  //                .readdata
		input  wire        node_131073_mem_write,     //                .write
		input  wire [15:0] node_131073_mem_writedata, //                .writedata
		input  wire [14:0] node_131074_mem_address,   // node_131074_mem.address
		output wire [15:0] node_131074_mem_readdata,  //                .readdata
		input  wire        node_131074_mem_write,     //                .write
		input  wire [15:0] node_131074_mem_writedata, //                .writedata
		input  wire [14:0] node_131075_mem_address,   // node_131075_mem.address
		output wire [15:0] node_131075_mem_readdata,  //                .readdata
		input  wire        node_131075_mem_write,     //                .write
		input  wire [15:0] node_131075_mem_writedata, //                .writedata
		input  wire [14:0] node_131076_mem_address,   // node_131076_mem.address
		output wire [15:0] node_131076_mem_readdata,  //                .readdata
		input  wire        node_131076_mem_write,     //                .write
		input  wire [15:0] node_131076_mem_writedata, //                .writedata
		input  wire [14:0] node_131077_mem_address,   // node_131077_mem.address
		output wire [15:0] node_131077_mem_readdata,  //                .readdata
		input  wire        node_131077_mem_write,     //                .write
		input  wire [15:0] node_131077_mem_writedata, //                .writedata
		input  wire [14:0] node_131078_mem_address,   // node_131078_mem.address
		output wire [15:0] node_131078_mem_readdata,  //                .readdata
		input  wire        node_131078_mem_write,     //                .write
		input  wire [15:0] node_131078_mem_writedata, //                .writedata
		input  wire [14:0] node_131079_mem_address,   // node_131079_mem.address
		output wire [15:0] node_131079_mem_readdata,  //                .readdata
		input  wire        node_131079_mem_write,     //                .write
		input  wire [15:0] node_131079_mem_writedata, //                .writedata
		input  wire [14:0] node_131080_mem_address,   // node_131080_mem.address
		output wire [15:0] node_131080_mem_readdata,  //                .readdata
		input  wire        node_131080_mem_write,     //                .write
		input  wire [15:0] node_131080_mem_writedata, //                .writedata
		input  wire [14:0] node_1_mem_address,        //      node_1_mem.address
		output wire [15:0] node_1_mem_readdata,       //                .readdata
		input  wire        node_1_mem_write,          //                .write
		input  wire [15:0] node_1_mem_writedata,      //                .writedata
		input  wire [14:0] node_2_mem_address,        //      node_2_mem.address
		output wire [15:0] node_2_mem_readdata,       //                .readdata
		input  wire        node_2_mem_write,          //                .write
		input  wire [15:0] node_2_mem_writedata,      //                .writedata
		input  wire [14:0] node_3_mem_address,        //      node_3_mem.address
		output wire [15:0] node_3_mem_readdata,       //                .readdata
		input  wire        node_3_mem_write,          //                .write
		input  wire [15:0] node_3_mem_writedata,      //                .writedata
		input  wire [14:0] node_4_mem_address,        //      node_4_mem.address
		output wire [15:0] node_4_mem_readdata,       //                .readdata
		input  wire        node_4_mem_write,          //                .write
		input  wire [15:0] node_4_mem_writedata,      //                .writedata
		input  wire [14:0] node_5_mem_address,        //      node_5_mem.address
		output wire [15:0] node_5_mem_readdata,       //                .readdata
		input  wire        node_5_mem_write,          //                .write
		input  wire [15:0] node_5_mem_writedata,      //                .writedata
		input  wire [14:0] node_65536_mem_address,    //  node_65536_mem.address
		output wire [15:0] node_65536_mem_readdata,   //                .readdata
		input  wire        node_65536_mem_write,      //                .write
		input  wire [15:0] node_65536_mem_writedata,  //                .writedata
		input  wire [14:0] node_65537_mem_address,    //  node_65537_mem.address
		output wire [15:0] node_65537_mem_readdata,   //                .readdata
		input  wire        node_65537_mem_write,      //                .write
		input  wire [15:0] node_65537_mem_writedata,  //                .writedata
		input  wire [14:0] node_65538_mem_address,    //  node_65538_mem.address
		output wire [15:0] node_65538_mem_readdata,   //                .readdata
		input  wire        node_65538_mem_write,      //                .write
		input  wire [15:0] node_65538_mem_writedata,  //                .writedata
		input  wire [14:0] node_65539_mem_address,    //  node_65539_mem.address
		output wire [15:0] node_65539_mem_readdata,   //                .readdata
		input  wire        node_65539_mem_write,      //                .write
		input  wire [15:0] node_65539_mem_writedata,  //                .writedata
		input  wire [14:0] node_65540_mem_address,    //  node_65540_mem.address
		output wire [15:0] node_65540_mem_readdata,   //                .readdata
		input  wire        node_65540_mem_write,      //                .write
		input  wire [15:0] node_65540_mem_writedata,  //                .writedata
		input  wire [14:0] node_65541_mem_address,    //  node_65541_mem.address
		output wire [15:0] node_65541_mem_readdata,   //                .readdata
		input  wire        node_65541_mem_write,      //                .write
		input  wire [15:0] node_65541_mem_writedata,  //                .writedata
		input  wire [14:0] node_65542_mem_address,    //  node_65542_mem.address
		output wire [15:0] node_65542_mem_readdata,   //                .readdata
		input  wire        node_65542_mem_write,      //                .write
		input  wire [15:0] node_65542_mem_writedata,  //                .writedata
		input  wire [14:0] node_65543_mem_address,    //  node_65543_mem.address
		output wire [15:0] node_65543_mem_readdata,   //                .readdata
		input  wire        node_65543_mem_write,      //                .write
		input  wire [15:0] node_65543_mem_writedata,  //                .writedata
		input  wire [14:0] node_65544_mem_address,    //  node_65544_mem.address
		output wire [15:0] node_65544_mem_readdata,   //                .readdata
		input  wire        node_65544_mem_write,      //                .write
		input  wire [15:0] node_65544_mem_writedata,  //                .writedata
		input  wire [14:0] node_6_mem_address,        //      node_6_mem.address
		output wire [15:0] node_6_mem_readdata,       //                .readdata
		input  wire        node_6_mem_write,          //                .write
		input  wire [15:0] node_6_mem_writedata,      //                .writedata
		input  wire [14:0] node_7_mem_address,        //      node_7_mem.address
		output wire [15:0] node_7_mem_readdata,       //                .readdata
		input  wire        node_7_mem_write,          //                .write
		input  wire [15:0] node_7_mem_writedata,      //                .writedata
		input  wire [14:0] node_8_mem_address,        //      node_8_mem.address
		output wire [15:0] node_8_mem_readdata,       //                .readdata
		input  wire        node_8_mem_write,          //                .write
		input  wire [15:0] node_8_mem_writedata,      //                .writedata
		input  wire        reset_reset_n,             //           reset.reset_n
		input  wire        reset_13_reset_n           //        reset_13.reset_n
	);

	wire         node_0_output_east_valid;               // node_0:output_east_valid -> node_1:input_west_valid
	wire  [31:0] node_0_output_east_data;                // node_0:output_east_data -> node_1:input_west_data
	wire         node_0_output_east_ready;               // node_1:input_west_ready -> node_0:output_east_ready
	wire         node_0_output_east_startofpacket;       // node_0:output_east_startofpacket -> node_1:input_west_startofpacket
	wire         node_0_output_east_endofpacket;         // node_0:output_east_endofpacket -> node_1:input_west_endofpacket
	wire   [1:0] node_0_output_east_empty;               // node_0:output_east_empty -> node_1:input_west_empty
	wire         node_1_output_east_valid;               // node_1:output_east_valid -> node_2:input_west_valid
	wire  [31:0] node_1_output_east_data;                // node_1:output_east_data -> node_2:input_west_data
	wire         node_1_output_east_ready;               // node_2:input_west_ready -> node_1:output_east_ready
	wire         node_1_output_east_startofpacket;       // node_1:output_east_startofpacket -> node_2:input_west_startofpacket
	wire         node_1_output_east_endofpacket;         // node_1:output_east_endofpacket -> node_2:input_west_endofpacket
	wire   [1:0] node_1_output_east_empty;               // node_1:output_east_empty -> node_2:input_west_empty
	wire         node_65536_output_east_valid;           // node_65536:output_east_valid -> node_65537:input_west_valid
	wire  [31:0] node_65536_output_east_data;            // node_65536:output_east_data -> node_65537:input_west_data
	wire         node_65536_output_east_ready;           // node_65537:input_west_ready -> node_65536:output_east_ready
	wire         node_65536_output_east_startofpacket;   // node_65536:output_east_startofpacket -> node_65537:input_west_startofpacket
	wire         node_65536_output_east_endofpacket;     // node_65536:output_east_endofpacket -> node_65537:input_west_endofpacket
	wire   [1:0] node_65536_output_east_empty;           // node_65536:output_east_empty -> node_65537:input_west_empty
	wire         node_65537_output_east_valid;           // node_65537:output_east_valid -> node_65538:input_west_valid
	wire  [31:0] node_65537_output_east_data;            // node_65537:output_east_data -> node_65538:input_west_data
	wire         node_65537_output_east_ready;           // node_65538:input_west_ready -> node_65537:output_east_ready
	wire         node_65537_output_east_startofpacket;   // node_65537:output_east_startofpacket -> node_65538:input_west_startofpacket
	wire         node_65537_output_east_endofpacket;     // node_65537:output_east_endofpacket -> node_65538:input_west_endofpacket
	wire   [1:0] node_65537_output_east_empty;           // node_65537:output_east_empty -> node_65538:input_west_empty
	wire         node_131072_output_east_valid;          // node_131072:output_east_valid -> node_131073:input_west_valid
	wire  [31:0] node_131072_output_east_data;           // node_131072:output_east_data -> node_131073:input_west_data
	wire         node_131072_output_east_ready;          // node_131073:input_west_ready -> node_131072:output_east_ready
	wire         node_131072_output_east_startofpacket;  // node_131072:output_east_startofpacket -> node_131073:input_west_startofpacket
	wire         node_131072_output_east_endofpacket;    // node_131072:output_east_endofpacket -> node_131073:input_west_endofpacket
	wire   [1:0] node_131072_output_east_empty;          // node_131072:output_east_empty -> node_131073:input_west_empty
	wire         node_131073_output_east_valid;          // node_131073:output_east_valid -> node_131074:input_west_valid
	wire  [31:0] node_131073_output_east_data;           // node_131073:output_east_data -> node_131074:input_west_data
	wire         node_131073_output_east_ready;          // node_131074:input_west_ready -> node_131073:output_east_ready
	wire         node_131073_output_east_startofpacket;  // node_131073:output_east_startofpacket -> node_131074:input_west_startofpacket
	wire         node_131073_output_east_endofpacket;    // node_131073:output_east_endofpacket -> node_131074:input_west_endofpacket
	wire   [1:0] node_131073_output_east_empty;          // node_131073:output_east_empty -> node_131074:input_west_empty
	wire         node_2_output_east_valid;               // node_2:output_east_valid -> node_3:input_west_valid
	wire  [31:0] node_2_output_east_data;                // node_2:output_east_data -> node_3:input_west_data
	wire         node_2_output_east_ready;               // node_3:input_west_ready -> node_2:output_east_ready
	wire         node_2_output_east_startofpacket;       // node_2:output_east_startofpacket -> node_3:input_west_startofpacket
	wire         node_2_output_east_endofpacket;         // node_2:output_east_endofpacket -> node_3:input_west_endofpacket
	wire   [1:0] node_2_output_east_empty;               // node_2:output_east_empty -> node_3:input_west_empty
	wire         node_3_output_east_valid;               // node_3:output_east_valid -> node_4:input_west_valid
	wire  [31:0] node_3_output_east_data;                // node_3:output_east_data -> node_4:input_west_data
	wire         node_3_output_east_ready;               // node_4:input_west_ready -> node_3:output_east_ready
	wire         node_3_output_east_startofpacket;       // node_3:output_east_startofpacket -> node_4:input_west_startofpacket
	wire         node_3_output_east_endofpacket;         // node_3:output_east_endofpacket -> node_4:input_west_endofpacket
	wire   [1:0] node_3_output_east_empty;               // node_3:output_east_empty -> node_4:input_west_empty
	wire         node_4_output_east_valid;               // node_4:output_east_valid -> node_5:input_west_valid
	wire  [31:0] node_4_output_east_data;                // node_4:output_east_data -> node_5:input_west_data
	wire         node_4_output_east_ready;               // node_5:input_west_ready -> node_4:output_east_ready
	wire         node_4_output_east_startofpacket;       // node_4:output_east_startofpacket -> node_5:input_west_startofpacket
	wire         node_4_output_east_endofpacket;         // node_4:output_east_endofpacket -> node_5:input_west_endofpacket
	wire   [1:0] node_4_output_east_empty;               // node_4:output_east_empty -> node_5:input_west_empty
	wire         node_5_output_east_valid;               // node_5:output_east_valid -> node_6:input_west_valid
	wire  [31:0] node_5_output_east_data;                // node_5:output_east_data -> node_6:input_west_data
	wire         node_5_output_east_ready;               // node_6:input_west_ready -> node_5:output_east_ready
	wire         node_5_output_east_startofpacket;       // node_5:output_east_startofpacket -> node_6:input_west_startofpacket
	wire         node_5_output_east_endofpacket;         // node_5:output_east_endofpacket -> node_6:input_west_endofpacket
	wire   [1:0] node_5_output_east_empty;               // node_5:output_east_empty -> node_6:input_west_empty
	wire         node_6_output_east_valid;               // node_6:output_east_valid -> node_7:input_west_valid
	wire  [31:0] node_6_output_east_data;                // node_6:output_east_data -> node_7:input_west_data
	wire         node_6_output_east_ready;               // node_7:input_west_ready -> node_6:output_east_ready
	wire         node_6_output_east_startofpacket;       // node_6:output_east_startofpacket -> node_7:input_west_startofpacket
	wire         node_6_output_east_endofpacket;         // node_6:output_east_endofpacket -> node_7:input_west_endofpacket
	wire   [1:0] node_6_output_east_empty;               // node_6:output_east_empty -> node_7:input_west_empty
	wire         node_7_output_east_valid;               // node_7:output_east_valid -> node_8:input_west_valid
	wire  [31:0] node_7_output_east_data;                // node_7:output_east_data -> node_8:input_west_data
	wire         node_7_output_east_ready;               // node_8:input_west_ready -> node_7:output_east_ready
	wire         node_7_output_east_startofpacket;       // node_7:output_east_startofpacket -> node_8:input_west_startofpacket
	wire         node_7_output_east_endofpacket;         // node_7:output_east_endofpacket -> node_8:input_west_endofpacket
	wire   [1:0] node_7_output_east_empty;               // node_7:output_east_empty -> node_8:input_west_empty
	wire         node_65538_output_east_valid;           // node_65538:output_east_valid -> node_65539:input_west_valid
	wire  [31:0] node_65538_output_east_data;            // node_65538:output_east_data -> node_65539:input_west_data
	wire         node_65538_output_east_ready;           // node_65539:input_west_ready -> node_65538:output_east_ready
	wire         node_65538_output_east_startofpacket;   // node_65538:output_east_startofpacket -> node_65539:input_west_startofpacket
	wire         node_65538_output_east_endofpacket;     // node_65538:output_east_endofpacket -> node_65539:input_west_endofpacket
	wire   [1:0] node_65538_output_east_empty;           // node_65538:output_east_empty -> node_65539:input_west_empty
	wire         node_65539_output_east_valid;           // node_65539:output_east_valid -> node_65540:input_west_valid
	wire  [31:0] node_65539_output_east_data;            // node_65539:output_east_data -> node_65540:input_west_data
	wire         node_65539_output_east_ready;           // node_65540:input_west_ready -> node_65539:output_east_ready
	wire         node_65539_output_east_startofpacket;   // node_65539:output_east_startofpacket -> node_65540:input_west_startofpacket
	wire         node_65539_output_east_endofpacket;     // node_65539:output_east_endofpacket -> node_65540:input_west_endofpacket
	wire   [1:0] node_65539_output_east_empty;           // node_65539:output_east_empty -> node_65540:input_west_empty
	wire         node_65540_output_east_valid;           // node_65540:output_east_valid -> node_65541:input_west_valid
	wire  [31:0] node_65540_output_east_data;            // node_65540:output_east_data -> node_65541:input_west_data
	wire         node_65540_output_east_ready;           // node_65541:input_west_ready -> node_65540:output_east_ready
	wire         node_65540_output_east_startofpacket;   // node_65540:output_east_startofpacket -> node_65541:input_west_startofpacket
	wire         node_65540_output_east_endofpacket;     // node_65540:output_east_endofpacket -> node_65541:input_west_endofpacket
	wire   [1:0] node_65540_output_east_empty;           // node_65540:output_east_empty -> node_65541:input_west_empty
	wire         node_65541_output_east_valid;           // node_65541:output_east_valid -> node_65542:input_west_valid
	wire  [31:0] node_65541_output_east_data;            // node_65541:output_east_data -> node_65542:input_west_data
	wire         node_65541_output_east_ready;           // node_65542:input_west_ready -> node_65541:output_east_ready
	wire         node_65541_output_east_startofpacket;   // node_65541:output_east_startofpacket -> node_65542:input_west_startofpacket
	wire         node_65541_output_east_endofpacket;     // node_65541:output_east_endofpacket -> node_65542:input_west_endofpacket
	wire   [1:0] node_65541_output_east_empty;           // node_65541:output_east_empty -> node_65542:input_west_empty
	wire         node_65542_output_east_valid;           // node_65542:output_east_valid -> node_65543:input_west_valid
	wire  [31:0] node_65542_output_east_data;            // node_65542:output_east_data -> node_65543:input_west_data
	wire         node_65542_output_east_ready;           // node_65543:input_west_ready -> node_65542:output_east_ready
	wire         node_65542_output_east_startofpacket;   // node_65542:output_east_startofpacket -> node_65543:input_west_startofpacket
	wire         node_65542_output_east_endofpacket;     // node_65542:output_east_endofpacket -> node_65543:input_west_endofpacket
	wire   [1:0] node_65542_output_east_empty;           // node_65542:output_east_empty -> node_65543:input_west_empty
	wire         node_65543_output_east_valid;           // node_65543:output_east_valid -> node_65544:input_west_valid
	wire  [31:0] node_65543_output_east_data;            // node_65543:output_east_data -> node_65544:input_west_data
	wire         node_65543_output_east_ready;           // node_65544:input_west_ready -> node_65543:output_east_ready
	wire         node_65543_output_east_startofpacket;   // node_65543:output_east_startofpacket -> node_65544:input_west_startofpacket
	wire         node_65543_output_east_endofpacket;     // node_65543:output_east_endofpacket -> node_65544:input_west_endofpacket
	wire   [1:0] node_65543_output_east_empty;           // node_65543:output_east_empty -> node_65544:input_west_empty
	wire         node_131074_output_east_valid;          // node_131074:output_east_valid -> node_131075:input_west_valid
	wire  [31:0] node_131074_output_east_data;           // node_131074:output_east_data -> node_131075:input_west_data
	wire         node_131074_output_east_ready;          // node_131075:input_west_ready -> node_131074:output_east_ready
	wire         node_131074_output_east_startofpacket;  // node_131074:output_east_startofpacket -> node_131075:input_west_startofpacket
	wire         node_131074_output_east_endofpacket;    // node_131074:output_east_endofpacket -> node_131075:input_west_endofpacket
	wire   [1:0] node_131074_output_east_empty;          // node_131074:output_east_empty -> node_131075:input_west_empty
	wire         node_131075_output_east_valid;          // node_131075:output_east_valid -> node_131076:input_west_valid
	wire  [31:0] node_131075_output_east_data;           // node_131075:output_east_data -> node_131076:input_west_data
	wire         node_131075_output_east_ready;          // node_131076:input_west_ready -> node_131075:output_east_ready
	wire         node_131075_output_east_startofpacket;  // node_131075:output_east_startofpacket -> node_131076:input_west_startofpacket
	wire         node_131075_output_east_endofpacket;    // node_131075:output_east_endofpacket -> node_131076:input_west_endofpacket
	wire   [1:0] node_131075_output_east_empty;          // node_131075:output_east_empty -> node_131076:input_west_empty
	wire         node_131076_output_east_valid;          // node_131076:output_east_valid -> node_131077:input_west_valid
	wire  [31:0] node_131076_output_east_data;           // node_131076:output_east_data -> node_131077:input_west_data
	wire         node_131076_output_east_ready;          // node_131077:input_west_ready -> node_131076:output_east_ready
	wire         node_131076_output_east_startofpacket;  // node_131076:output_east_startofpacket -> node_131077:input_west_startofpacket
	wire         node_131076_output_east_endofpacket;    // node_131076:output_east_endofpacket -> node_131077:input_west_endofpacket
	wire   [1:0] node_131076_output_east_empty;          // node_131076:output_east_empty -> node_131077:input_west_empty
	wire         node_131077_output_east_valid;          // node_131077:output_east_valid -> node_131078:input_west_valid
	wire  [31:0] node_131077_output_east_data;           // node_131077:output_east_data -> node_131078:input_west_data
	wire         node_131077_output_east_ready;          // node_131078:input_west_ready -> node_131077:output_east_ready
	wire         node_131077_output_east_startofpacket;  // node_131077:output_east_startofpacket -> node_131078:input_west_startofpacket
	wire         node_131077_output_east_endofpacket;    // node_131077:output_east_endofpacket -> node_131078:input_west_endofpacket
	wire   [1:0] node_131077_output_east_empty;          // node_131077:output_east_empty -> node_131078:input_west_empty
	wire         node_131079_output_east_valid;          // node_131079:output_east_valid -> node_131080:input_west_valid
	wire  [31:0] node_131079_output_east_data;           // node_131079:output_east_data -> node_131080:input_west_data
	wire         node_131079_output_east_ready;          // node_131080:input_west_ready -> node_131079:output_east_ready
	wire         node_131079_output_east_startofpacket;  // node_131079:output_east_startofpacket -> node_131080:input_west_startofpacket
	wire         node_131079_output_east_endofpacket;    // node_131079:output_east_endofpacket -> node_131080:input_west_endofpacket
	wire   [1:0] node_131079_output_east_empty;          // node_131079:output_east_empty -> node_131080:input_west_empty
	wire         node_131078_output_east_valid;          // node_131078:output_east_valid -> node_131079:input_west_valid
	wire  [31:0] node_131078_output_east_data;           // node_131078:output_east_data -> node_131079:input_west_data
	wire         node_131078_output_east_ready;          // node_131079:input_west_ready -> node_131078:output_east_ready
	wire         node_131078_output_east_startofpacket;  // node_131078:output_east_startofpacket -> node_131079:input_west_startofpacket
	wire         node_131078_output_east_endofpacket;    // node_131078:output_east_endofpacket -> node_131079:input_west_endofpacket
	wire   [1:0] node_131078_output_east_empty;          // node_131078:output_east_empty -> node_131079:input_west_empty
	wire         node_8_output_east_valid;               // node_8:output_east_valid -> terminal_east_0:valid
	wire  [31:0] node_8_output_east_data;                // node_8:output_east_data -> terminal_east_0:data
	wire         node_8_output_east_ready;               // terminal_east_0:ready -> node_8:output_east_ready
	wire         node_8_output_east_startofpacket;       // node_8:output_east_startofpacket -> terminal_east_0:startofpacket
	wire         node_8_output_east_endofpacket;         // node_8:output_east_endofpacket -> terminal_east_0:endofpacket
	wire   [1:0] node_8_output_east_empty;               // node_8:output_east_empty -> terminal_east_0:empty
	wire         node_131080_output_east_valid;          // node_131080:output_east_valid -> terminal_east_2:valid
	wire  [31:0] node_131080_output_east_data;           // node_131080:output_east_data -> terminal_east_2:data
	wire         node_131080_output_east_ready;          // terminal_east_2:ready -> node_131080:output_east_ready
	wire         node_131080_output_east_startofpacket;  // node_131080:output_east_startofpacket -> terminal_east_2:startofpacket
	wire         node_131080_output_east_endofpacket;    // node_131080:output_east_endofpacket -> terminal_east_2:endofpacket
	wire   [1:0] node_131080_output_east_empty;          // node_131080:output_east_empty -> terminal_east_2:empty
	wire         node_65544_output_east_valid;           // node_65544:output_east_valid -> terminal_east_1:valid
	wire  [31:0] node_65544_output_east_data;            // node_65544:output_east_data -> terminal_east_1:data
	wire         node_65544_output_east_ready;           // terminal_east_1:ready -> node_65544:output_east_ready
	wire         node_65544_output_east_startofpacket;   // node_65544:output_east_startofpacket -> terminal_east_1:startofpacket
	wire         node_65544_output_east_endofpacket;     // node_65544:output_east_endofpacket -> terminal_east_1:endofpacket
	wire   [1:0] node_65544_output_east_empty;           // node_65544:output_east_empty -> terminal_east_1:empty
	wire         node_65536_output_north_valid;          // node_65536:output_north_valid -> node_0:input_south_valid
	wire  [31:0] node_65536_output_north_data;           // node_65536:output_north_data -> node_0:input_south_data
	wire         node_65536_output_north_ready;          // node_0:input_south_ready -> node_65536:output_north_ready
	wire         node_65536_output_north_startofpacket;  // node_65536:output_north_startofpacket -> node_0:input_south_startofpacket
	wire         node_65536_output_north_endofpacket;    // node_65536:output_north_endofpacket -> node_0:input_south_endofpacket
	wire   [1:0] node_65536_output_north_empty;          // node_65536:output_north_empty -> node_0:input_south_empty
	wire         node_65537_output_north_valid;          // node_65537:output_north_valid -> node_1:input_south_valid
	wire  [31:0] node_65537_output_north_data;           // node_65537:output_north_data -> node_1:input_south_data
	wire         node_65537_output_north_ready;          // node_1:input_south_ready -> node_65537:output_north_ready
	wire         node_65537_output_north_startofpacket;  // node_65537:output_north_startofpacket -> node_1:input_south_startofpacket
	wire         node_65537_output_north_endofpacket;    // node_65537:output_north_endofpacket -> node_1:input_south_endofpacket
	wire   [1:0] node_65537_output_north_empty;          // node_65537:output_north_empty -> node_1:input_south_empty
	wire         node_65538_output_north_valid;          // node_65538:output_north_valid -> node_2:input_south_valid
	wire  [31:0] node_65538_output_north_data;           // node_65538:output_north_data -> node_2:input_south_data
	wire         node_65538_output_north_ready;          // node_2:input_south_ready -> node_65538:output_north_ready
	wire         node_65538_output_north_startofpacket;  // node_65538:output_north_startofpacket -> node_2:input_south_startofpacket
	wire         node_65538_output_north_endofpacket;    // node_65538:output_north_endofpacket -> node_2:input_south_endofpacket
	wire   [1:0] node_65538_output_north_empty;          // node_65538:output_north_empty -> node_2:input_south_empty
	wire         node_65539_output_north_valid;          // node_65539:output_north_valid -> node_3:input_south_valid
	wire  [31:0] node_65539_output_north_data;           // node_65539:output_north_data -> node_3:input_south_data
	wire         node_65539_output_north_ready;          // node_3:input_south_ready -> node_65539:output_north_ready
	wire         node_65539_output_north_startofpacket;  // node_65539:output_north_startofpacket -> node_3:input_south_startofpacket
	wire         node_65539_output_north_endofpacket;    // node_65539:output_north_endofpacket -> node_3:input_south_endofpacket
	wire   [1:0] node_65539_output_north_empty;          // node_65539:output_north_empty -> node_3:input_south_empty
	wire         node_65540_output_north_valid;          // node_65540:output_north_valid -> node_4:input_south_valid
	wire  [31:0] node_65540_output_north_data;           // node_65540:output_north_data -> node_4:input_south_data
	wire         node_65540_output_north_ready;          // node_4:input_south_ready -> node_65540:output_north_ready
	wire         node_65540_output_north_startofpacket;  // node_65540:output_north_startofpacket -> node_4:input_south_startofpacket
	wire         node_65540_output_north_endofpacket;    // node_65540:output_north_endofpacket -> node_4:input_south_endofpacket
	wire   [1:0] node_65540_output_north_empty;          // node_65540:output_north_empty -> node_4:input_south_empty
	wire         node_65541_output_north_valid;          // node_65541:output_north_valid -> node_5:input_south_valid
	wire  [31:0] node_65541_output_north_data;           // node_65541:output_north_data -> node_5:input_south_data
	wire         node_65541_output_north_ready;          // node_5:input_south_ready -> node_65541:output_north_ready
	wire         node_65541_output_north_startofpacket;  // node_65541:output_north_startofpacket -> node_5:input_south_startofpacket
	wire         node_65541_output_north_endofpacket;    // node_65541:output_north_endofpacket -> node_5:input_south_endofpacket
	wire   [1:0] node_65541_output_north_empty;          // node_65541:output_north_empty -> node_5:input_south_empty
	wire         node_65542_output_north_valid;          // node_65542:output_north_valid -> node_6:input_south_valid
	wire  [31:0] node_65542_output_north_data;           // node_65542:output_north_data -> node_6:input_south_data
	wire         node_65542_output_north_ready;          // node_6:input_south_ready -> node_65542:output_north_ready
	wire         node_65542_output_north_startofpacket;  // node_65542:output_north_startofpacket -> node_6:input_south_startofpacket
	wire         node_65542_output_north_endofpacket;    // node_65542:output_north_endofpacket -> node_6:input_south_endofpacket
	wire   [1:0] node_65542_output_north_empty;          // node_65542:output_north_empty -> node_6:input_south_empty
	wire         node_65543_output_north_valid;          // node_65543:output_north_valid -> node_7:input_south_valid
	wire  [31:0] node_65543_output_north_data;           // node_65543:output_north_data -> node_7:input_south_data
	wire         node_65543_output_north_ready;          // node_7:input_south_ready -> node_65543:output_north_ready
	wire         node_65543_output_north_startofpacket;  // node_65543:output_north_startofpacket -> node_7:input_south_startofpacket
	wire         node_65543_output_north_endofpacket;    // node_65543:output_north_endofpacket -> node_7:input_south_endofpacket
	wire   [1:0] node_65543_output_north_empty;          // node_65543:output_north_empty -> node_7:input_south_empty
	wire         node_65544_output_north_valid;          // node_65544:output_north_valid -> node_8:input_south_valid
	wire  [31:0] node_65544_output_north_data;           // node_65544:output_north_data -> node_8:input_south_data
	wire         node_65544_output_north_ready;          // node_8:input_south_ready -> node_65544:output_north_ready
	wire         node_65544_output_north_startofpacket;  // node_65544:output_north_startofpacket -> node_8:input_south_startofpacket
	wire         node_65544_output_north_endofpacket;    // node_65544:output_north_endofpacket -> node_8:input_south_endofpacket
	wire   [1:0] node_65544_output_north_empty;          // node_65544:output_north_empty -> node_8:input_south_empty
	wire         node_131072_output_north_valid;         // node_131072:output_north_valid -> node_65536:input_south_valid
	wire  [31:0] node_131072_output_north_data;          // node_131072:output_north_data -> node_65536:input_south_data
	wire         node_131072_output_north_ready;         // node_65536:input_south_ready -> node_131072:output_north_ready
	wire         node_131072_output_north_startofpacket; // node_131072:output_north_startofpacket -> node_65536:input_south_startofpacket
	wire         node_131072_output_north_endofpacket;   // node_131072:output_north_endofpacket -> node_65536:input_south_endofpacket
	wire   [1:0] node_131072_output_north_empty;         // node_131072:output_north_empty -> node_65536:input_south_empty
	wire         node_131073_output_north_valid;         // node_131073:output_north_valid -> node_65537:input_south_valid
	wire  [31:0] node_131073_output_north_data;          // node_131073:output_north_data -> node_65537:input_south_data
	wire         node_131073_output_north_ready;         // node_65537:input_south_ready -> node_131073:output_north_ready
	wire         node_131073_output_north_startofpacket; // node_131073:output_north_startofpacket -> node_65537:input_south_startofpacket
	wire         node_131073_output_north_endofpacket;   // node_131073:output_north_endofpacket -> node_65537:input_south_endofpacket
	wire   [1:0] node_131073_output_north_empty;         // node_131073:output_north_empty -> node_65537:input_south_empty
	wire         node_131074_output_north_valid;         // node_131074:output_north_valid -> node_65538:input_south_valid
	wire  [31:0] node_131074_output_north_data;          // node_131074:output_north_data -> node_65538:input_south_data
	wire         node_131074_output_north_ready;         // node_65538:input_south_ready -> node_131074:output_north_ready
	wire         node_131074_output_north_startofpacket; // node_131074:output_north_startofpacket -> node_65538:input_south_startofpacket
	wire         node_131074_output_north_endofpacket;   // node_131074:output_north_endofpacket -> node_65538:input_south_endofpacket
	wire   [1:0] node_131074_output_north_empty;         // node_131074:output_north_empty -> node_65538:input_south_empty
	wire         node_131075_output_north_valid;         // node_131075:output_north_valid -> node_65539:input_south_valid
	wire  [31:0] node_131075_output_north_data;          // node_131075:output_north_data -> node_65539:input_south_data
	wire         node_131075_output_north_ready;         // node_65539:input_south_ready -> node_131075:output_north_ready
	wire         node_131075_output_north_startofpacket; // node_131075:output_north_startofpacket -> node_65539:input_south_startofpacket
	wire         node_131075_output_north_endofpacket;   // node_131075:output_north_endofpacket -> node_65539:input_south_endofpacket
	wire   [1:0] node_131075_output_north_empty;         // node_131075:output_north_empty -> node_65539:input_south_empty
	wire         node_131076_output_north_valid;         // node_131076:output_north_valid -> node_65540:input_south_valid
	wire  [31:0] node_131076_output_north_data;          // node_131076:output_north_data -> node_65540:input_south_data
	wire         node_131076_output_north_ready;         // node_65540:input_south_ready -> node_131076:output_north_ready
	wire         node_131076_output_north_startofpacket; // node_131076:output_north_startofpacket -> node_65540:input_south_startofpacket
	wire         node_131076_output_north_endofpacket;   // node_131076:output_north_endofpacket -> node_65540:input_south_endofpacket
	wire   [1:0] node_131076_output_north_empty;         // node_131076:output_north_empty -> node_65540:input_south_empty
	wire         node_131077_output_north_valid;         // node_131077:output_north_valid -> node_65541:input_south_valid
	wire  [31:0] node_131077_output_north_data;          // node_131077:output_north_data -> node_65541:input_south_data
	wire         node_131077_output_north_ready;         // node_65541:input_south_ready -> node_131077:output_north_ready
	wire         node_131077_output_north_startofpacket; // node_131077:output_north_startofpacket -> node_65541:input_south_startofpacket
	wire         node_131077_output_north_endofpacket;   // node_131077:output_north_endofpacket -> node_65541:input_south_endofpacket
	wire   [1:0] node_131077_output_north_empty;         // node_131077:output_north_empty -> node_65541:input_south_empty
	wire         node_131078_output_north_valid;         // node_131078:output_north_valid -> node_65542:input_south_valid
	wire  [31:0] node_131078_output_north_data;          // node_131078:output_north_data -> node_65542:input_south_data
	wire         node_131078_output_north_ready;         // node_65542:input_south_ready -> node_131078:output_north_ready
	wire         node_131078_output_north_startofpacket; // node_131078:output_north_startofpacket -> node_65542:input_south_startofpacket
	wire         node_131078_output_north_endofpacket;   // node_131078:output_north_endofpacket -> node_65542:input_south_endofpacket
	wire   [1:0] node_131078_output_north_empty;         // node_131078:output_north_empty -> node_65542:input_south_empty
	wire         node_131079_output_north_valid;         // node_131079:output_north_valid -> node_65543:input_south_valid
	wire  [31:0] node_131079_output_north_data;          // node_131079:output_north_data -> node_65543:input_south_data
	wire         node_131079_output_north_ready;         // node_65543:input_south_ready -> node_131079:output_north_ready
	wire         node_131079_output_north_startofpacket; // node_131079:output_north_startofpacket -> node_65543:input_south_startofpacket
	wire         node_131079_output_north_endofpacket;   // node_131079:output_north_endofpacket -> node_65543:input_south_endofpacket
	wire   [1:0] node_131079_output_north_empty;         // node_131079:output_north_empty -> node_65543:input_south_empty
	wire         node_131080_output_north_valid;         // node_131080:output_north_valid -> node_65544:input_south_valid
	wire  [31:0] node_131080_output_north_data;          // node_131080:output_north_data -> node_65544:input_south_data
	wire         node_131080_output_north_ready;         // node_65544:input_south_ready -> node_131080:output_north_ready
	wire         node_131080_output_north_startofpacket; // node_131080:output_north_startofpacket -> node_65544:input_south_startofpacket
	wire         node_131080_output_north_endofpacket;   // node_131080:output_north_endofpacket -> node_65544:input_south_endofpacket
	wire   [1:0] node_131080_output_north_empty;         // node_131080:output_north_empty -> node_65544:input_south_empty
	wire         node_0_output_north_valid;              // node_0:output_north_valid -> terminal_north_0:valid
	wire  [31:0] node_0_output_north_data;               // node_0:output_north_data -> terminal_north_0:data
	wire         node_0_output_north_ready;              // terminal_north_0:ready -> node_0:output_north_ready
	wire         node_0_output_north_startofpacket;      // node_0:output_north_startofpacket -> terminal_north_0:startofpacket
	wire         node_0_output_north_endofpacket;        // node_0:output_north_endofpacket -> terminal_north_0:endofpacket
	wire   [1:0] node_0_output_north_empty;              // node_0:output_north_empty -> terminal_north_0:empty
	wire         node_1_output_north_valid;              // node_1:output_north_valid -> terminal_north_1:valid
	wire  [31:0] node_1_output_north_data;               // node_1:output_north_data -> terminal_north_1:data
	wire         node_1_output_north_ready;              // terminal_north_1:ready -> node_1:output_north_ready
	wire         node_1_output_north_startofpacket;      // node_1:output_north_startofpacket -> terminal_north_1:startofpacket
	wire         node_1_output_north_endofpacket;        // node_1:output_north_endofpacket -> terminal_north_1:endofpacket
	wire   [1:0] node_1_output_north_empty;              // node_1:output_north_empty -> terminal_north_1:empty
	wire         node_2_output_north_valid;              // node_2:output_north_valid -> terminal_north_2:valid
	wire  [31:0] node_2_output_north_data;               // node_2:output_north_data -> terminal_north_2:data
	wire         node_2_output_north_ready;              // terminal_north_2:ready -> node_2:output_north_ready
	wire         node_2_output_north_startofpacket;      // node_2:output_north_startofpacket -> terminal_north_2:startofpacket
	wire         node_2_output_north_endofpacket;        // node_2:output_north_endofpacket -> terminal_north_2:endofpacket
	wire   [1:0] node_2_output_north_empty;              // node_2:output_north_empty -> terminal_north_2:empty
	wire         node_3_output_north_valid;              // node_3:output_north_valid -> terminal_north_3:valid
	wire  [31:0] node_3_output_north_data;               // node_3:output_north_data -> terminal_north_3:data
	wire         node_3_output_north_ready;              // terminal_north_3:ready -> node_3:output_north_ready
	wire         node_3_output_north_startofpacket;      // node_3:output_north_startofpacket -> terminal_north_3:startofpacket
	wire         node_3_output_north_endofpacket;        // node_3:output_north_endofpacket -> terminal_north_3:endofpacket
	wire   [1:0] node_3_output_north_empty;              // node_3:output_north_empty -> terminal_north_3:empty
	wire         node_4_output_north_valid;              // node_4:output_north_valid -> terminal_north_4:valid
	wire  [31:0] node_4_output_north_data;               // node_4:output_north_data -> terminal_north_4:data
	wire         node_4_output_north_ready;              // terminal_north_4:ready -> node_4:output_north_ready
	wire         node_4_output_north_startofpacket;      // node_4:output_north_startofpacket -> terminal_north_4:startofpacket
	wire         node_4_output_north_endofpacket;        // node_4:output_north_endofpacket -> terminal_north_4:endofpacket
	wire   [1:0] node_4_output_north_empty;              // node_4:output_north_empty -> terminal_north_4:empty
	wire         node_5_output_north_valid;              // node_5:output_north_valid -> terminal_north_5:valid
	wire  [31:0] node_5_output_north_data;               // node_5:output_north_data -> terminal_north_5:data
	wire         node_5_output_north_ready;              // terminal_north_5:ready -> node_5:output_north_ready
	wire         node_5_output_north_startofpacket;      // node_5:output_north_startofpacket -> terminal_north_5:startofpacket
	wire         node_5_output_north_endofpacket;        // node_5:output_north_endofpacket -> terminal_north_5:endofpacket
	wire   [1:0] node_5_output_north_empty;              // node_5:output_north_empty -> terminal_north_5:empty
	wire         node_6_output_north_valid;              // node_6:output_north_valid -> terminal_north_6:valid
	wire  [31:0] node_6_output_north_data;               // node_6:output_north_data -> terminal_north_6:data
	wire         node_6_output_north_ready;              // terminal_north_6:ready -> node_6:output_north_ready
	wire         node_6_output_north_startofpacket;      // node_6:output_north_startofpacket -> terminal_north_6:startofpacket
	wire         node_6_output_north_endofpacket;        // node_6:output_north_endofpacket -> terminal_north_6:endofpacket
	wire   [1:0] node_6_output_north_empty;              // node_6:output_north_empty -> terminal_north_6:empty
	wire         node_7_output_north_valid;              // node_7:output_north_valid -> terminal_north_7:valid
	wire  [31:0] node_7_output_north_data;               // node_7:output_north_data -> terminal_north_7:data
	wire         node_7_output_north_ready;              // terminal_north_7:ready -> node_7:output_north_ready
	wire         node_7_output_north_startofpacket;      // node_7:output_north_startofpacket -> terminal_north_7:startofpacket
	wire         node_7_output_north_endofpacket;        // node_7:output_north_endofpacket -> terminal_north_7:endofpacket
	wire   [1:0] node_7_output_north_empty;              // node_7:output_north_empty -> terminal_north_7:empty
	wire         node_8_output_north_valid;              // node_8:output_north_valid -> terminal_north_8:valid
	wire  [31:0] node_8_output_north_data;               // node_8:output_north_data -> terminal_north_8:data
	wire         node_8_output_north_ready;              // terminal_north_8:ready -> node_8:output_north_ready
	wire         node_8_output_north_startofpacket;      // node_8:output_north_startofpacket -> terminal_north_8:startofpacket
	wire         node_8_output_north_endofpacket;        // node_8:output_north_endofpacket -> terminal_north_8:endofpacket
	wire   [1:0] node_8_output_north_empty;              // node_8:output_north_empty -> terminal_north_8:empty
	wire         node_0_output_south_valid;              // node_0:output_south_valid -> node_65536:input_north_valid
	wire  [31:0] node_0_output_south_data;               // node_0:output_south_data -> node_65536:input_north_data
	wire         node_0_output_south_ready;              // node_65536:input_north_ready -> node_0:output_south_ready
	wire         node_0_output_south_startofpacket;      // node_0:output_south_startofpacket -> node_65536:input_north_startofpacket
	wire         node_0_output_south_endofpacket;        // node_0:output_south_endofpacket -> node_65536:input_north_endofpacket
	wire   [1:0] node_0_output_south_empty;              // node_0:output_south_empty -> node_65536:input_north_empty
	wire         node_1_output_south_valid;              // node_1:output_south_valid -> node_65537:input_north_valid
	wire  [31:0] node_1_output_south_data;               // node_1:output_south_data -> node_65537:input_north_data
	wire         node_1_output_south_ready;              // node_65537:input_north_ready -> node_1:output_south_ready
	wire         node_1_output_south_startofpacket;      // node_1:output_south_startofpacket -> node_65537:input_north_startofpacket
	wire         node_1_output_south_endofpacket;        // node_1:output_south_endofpacket -> node_65537:input_north_endofpacket
	wire   [1:0] node_1_output_south_empty;              // node_1:output_south_empty -> node_65537:input_north_empty
	wire         node_2_output_south_valid;              // node_2:output_south_valid -> node_65538:input_north_valid
	wire  [31:0] node_2_output_south_data;               // node_2:output_south_data -> node_65538:input_north_data
	wire         node_2_output_south_ready;              // node_65538:input_north_ready -> node_2:output_south_ready
	wire         node_2_output_south_startofpacket;      // node_2:output_south_startofpacket -> node_65538:input_north_startofpacket
	wire         node_2_output_south_endofpacket;        // node_2:output_south_endofpacket -> node_65538:input_north_endofpacket
	wire   [1:0] node_2_output_south_empty;              // node_2:output_south_empty -> node_65538:input_north_empty
	wire         node_65536_output_south_valid;          // node_65536:output_south_valid -> node_131072:input_north_valid
	wire  [31:0] node_65536_output_south_data;           // node_65536:output_south_data -> node_131072:input_north_data
	wire         node_65536_output_south_ready;          // node_131072:input_north_ready -> node_65536:output_south_ready
	wire         node_65536_output_south_startofpacket;  // node_65536:output_south_startofpacket -> node_131072:input_north_startofpacket
	wire         node_65536_output_south_endofpacket;    // node_65536:output_south_endofpacket -> node_131072:input_north_endofpacket
	wire   [1:0] node_65536_output_south_empty;          // node_65536:output_south_empty -> node_131072:input_north_empty
	wire         node_65537_output_south_valid;          // node_65537:output_south_valid -> node_131073:input_north_valid
	wire  [31:0] node_65537_output_south_data;           // node_65537:output_south_data -> node_131073:input_north_data
	wire         node_65537_output_south_ready;          // node_131073:input_north_ready -> node_65537:output_south_ready
	wire         node_65537_output_south_startofpacket;  // node_65537:output_south_startofpacket -> node_131073:input_north_startofpacket
	wire         node_65537_output_south_endofpacket;    // node_65537:output_south_endofpacket -> node_131073:input_north_endofpacket
	wire   [1:0] node_65537_output_south_empty;          // node_65537:output_south_empty -> node_131073:input_north_empty
	wire         node_65538_output_south_valid;          // node_65538:output_south_valid -> node_131074:input_north_valid
	wire  [31:0] node_65538_output_south_data;           // node_65538:output_south_data -> node_131074:input_north_data
	wire         node_65538_output_south_ready;          // node_131074:input_north_ready -> node_65538:output_south_ready
	wire         node_65538_output_south_startofpacket;  // node_65538:output_south_startofpacket -> node_131074:input_north_startofpacket
	wire         node_65538_output_south_endofpacket;    // node_65538:output_south_endofpacket -> node_131074:input_north_endofpacket
	wire   [1:0] node_65538_output_south_empty;          // node_65538:output_south_empty -> node_131074:input_north_empty
	wire         node_3_output_south_valid;              // node_3:output_south_valid -> node_65539:input_north_valid
	wire  [31:0] node_3_output_south_data;               // node_3:output_south_data -> node_65539:input_north_data
	wire         node_3_output_south_ready;              // node_65539:input_north_ready -> node_3:output_south_ready
	wire         node_3_output_south_startofpacket;      // node_3:output_south_startofpacket -> node_65539:input_north_startofpacket
	wire         node_3_output_south_endofpacket;        // node_3:output_south_endofpacket -> node_65539:input_north_endofpacket
	wire   [1:0] node_3_output_south_empty;              // node_3:output_south_empty -> node_65539:input_north_empty
	wire         node_4_output_south_valid;              // node_4:output_south_valid -> node_65540:input_north_valid
	wire  [31:0] node_4_output_south_data;               // node_4:output_south_data -> node_65540:input_north_data
	wire         node_4_output_south_ready;              // node_65540:input_north_ready -> node_4:output_south_ready
	wire         node_4_output_south_startofpacket;      // node_4:output_south_startofpacket -> node_65540:input_north_startofpacket
	wire         node_4_output_south_endofpacket;        // node_4:output_south_endofpacket -> node_65540:input_north_endofpacket
	wire   [1:0] node_4_output_south_empty;              // node_4:output_south_empty -> node_65540:input_north_empty
	wire         node_5_output_south_valid;              // node_5:output_south_valid -> node_65541:input_north_valid
	wire  [31:0] node_5_output_south_data;               // node_5:output_south_data -> node_65541:input_north_data
	wire         node_5_output_south_ready;              // node_65541:input_north_ready -> node_5:output_south_ready
	wire         node_5_output_south_startofpacket;      // node_5:output_south_startofpacket -> node_65541:input_north_startofpacket
	wire         node_5_output_south_endofpacket;        // node_5:output_south_endofpacket -> node_65541:input_north_endofpacket
	wire   [1:0] node_5_output_south_empty;              // node_5:output_south_empty -> node_65541:input_north_empty
	wire         node_6_output_south_valid;              // node_6:output_south_valid -> node_65542:input_north_valid
	wire  [31:0] node_6_output_south_data;               // node_6:output_south_data -> node_65542:input_north_data
	wire         node_6_output_south_ready;              // node_65542:input_north_ready -> node_6:output_south_ready
	wire         node_6_output_south_startofpacket;      // node_6:output_south_startofpacket -> node_65542:input_north_startofpacket
	wire         node_6_output_south_endofpacket;        // node_6:output_south_endofpacket -> node_65542:input_north_endofpacket
	wire   [1:0] node_6_output_south_empty;              // node_6:output_south_empty -> node_65542:input_north_empty
	wire         node_7_output_south_valid;              // node_7:output_south_valid -> node_65543:input_north_valid
	wire  [31:0] node_7_output_south_data;               // node_7:output_south_data -> node_65543:input_north_data
	wire         node_7_output_south_ready;              // node_65543:input_north_ready -> node_7:output_south_ready
	wire         node_7_output_south_startofpacket;      // node_7:output_south_startofpacket -> node_65543:input_north_startofpacket
	wire         node_7_output_south_endofpacket;        // node_7:output_south_endofpacket -> node_65543:input_north_endofpacket
	wire   [1:0] node_7_output_south_empty;              // node_7:output_south_empty -> node_65543:input_north_empty
	wire         node_8_output_south_valid;              // node_8:output_south_valid -> node_65544:input_north_valid
	wire  [31:0] node_8_output_south_data;               // node_8:output_south_data -> node_65544:input_north_data
	wire         node_8_output_south_ready;              // node_65544:input_north_ready -> node_8:output_south_ready
	wire         node_8_output_south_startofpacket;      // node_8:output_south_startofpacket -> node_65544:input_north_startofpacket
	wire         node_8_output_south_endofpacket;        // node_8:output_south_endofpacket -> node_65544:input_north_endofpacket
	wire   [1:0] node_8_output_south_empty;              // node_8:output_south_empty -> node_65544:input_north_empty
	wire         node_65539_output_south_valid;          // node_65539:output_south_valid -> node_131075:input_north_valid
	wire  [31:0] node_65539_output_south_data;           // node_65539:output_south_data -> node_131075:input_north_data
	wire         node_65539_output_south_ready;          // node_131075:input_north_ready -> node_65539:output_south_ready
	wire         node_65539_output_south_startofpacket;  // node_65539:output_south_startofpacket -> node_131075:input_north_startofpacket
	wire         node_65539_output_south_endofpacket;    // node_65539:output_south_endofpacket -> node_131075:input_north_endofpacket
	wire   [1:0] node_65539_output_south_empty;          // node_65539:output_south_empty -> node_131075:input_north_empty
	wire         node_65540_output_south_valid;          // node_65540:output_south_valid -> node_131076:input_north_valid
	wire  [31:0] node_65540_output_south_data;           // node_65540:output_south_data -> node_131076:input_north_data
	wire         node_65540_output_south_ready;          // node_131076:input_north_ready -> node_65540:output_south_ready
	wire         node_65540_output_south_startofpacket;  // node_65540:output_south_startofpacket -> node_131076:input_north_startofpacket
	wire         node_65540_output_south_endofpacket;    // node_65540:output_south_endofpacket -> node_131076:input_north_endofpacket
	wire   [1:0] node_65540_output_south_empty;          // node_65540:output_south_empty -> node_131076:input_north_empty
	wire         node_65541_output_south_valid;          // node_65541:output_south_valid -> node_131077:input_north_valid
	wire  [31:0] node_65541_output_south_data;           // node_65541:output_south_data -> node_131077:input_north_data
	wire         node_65541_output_south_ready;          // node_131077:input_north_ready -> node_65541:output_south_ready
	wire         node_65541_output_south_startofpacket;  // node_65541:output_south_startofpacket -> node_131077:input_north_startofpacket
	wire         node_65541_output_south_endofpacket;    // node_65541:output_south_endofpacket -> node_131077:input_north_endofpacket
	wire   [1:0] node_65541_output_south_empty;          // node_65541:output_south_empty -> node_131077:input_north_empty
	wire         node_65542_output_south_valid;          // node_65542:output_south_valid -> node_131078:input_north_valid
	wire  [31:0] node_65542_output_south_data;           // node_65542:output_south_data -> node_131078:input_north_data
	wire         node_65542_output_south_ready;          // node_131078:input_north_ready -> node_65542:output_south_ready
	wire         node_65542_output_south_startofpacket;  // node_65542:output_south_startofpacket -> node_131078:input_north_startofpacket
	wire         node_65542_output_south_endofpacket;    // node_65542:output_south_endofpacket -> node_131078:input_north_endofpacket
	wire   [1:0] node_65542_output_south_empty;          // node_65542:output_south_empty -> node_131078:input_north_empty
	wire         node_65543_output_south_valid;          // node_65543:output_south_valid -> node_131079:input_north_valid
	wire  [31:0] node_65543_output_south_data;           // node_65543:output_south_data -> node_131079:input_north_data
	wire         node_65543_output_south_ready;          // node_131079:input_north_ready -> node_65543:output_south_ready
	wire         node_65543_output_south_startofpacket;  // node_65543:output_south_startofpacket -> node_131079:input_north_startofpacket
	wire         node_65543_output_south_endofpacket;    // node_65543:output_south_endofpacket -> node_131079:input_north_endofpacket
	wire   [1:0] node_65543_output_south_empty;          // node_65543:output_south_empty -> node_131079:input_north_empty
	wire         node_65544_output_south_valid;          // node_65544:output_south_valid -> node_131080:input_north_valid
	wire  [31:0] node_65544_output_south_data;           // node_65544:output_south_data -> node_131080:input_north_data
	wire         node_65544_output_south_ready;          // node_131080:input_north_ready -> node_65544:output_south_ready
	wire         node_65544_output_south_startofpacket;  // node_65544:output_south_startofpacket -> node_131080:input_north_startofpacket
	wire         node_65544_output_south_endofpacket;    // node_65544:output_south_endofpacket -> node_131080:input_north_endofpacket
	wire   [1:0] node_65544_output_south_empty;          // node_65544:output_south_empty -> node_131080:input_north_empty
	wire         node_131072_output_south_valid;         // node_131072:output_south_valid -> terminal_south_0:valid
	wire  [31:0] node_131072_output_south_data;          // node_131072:output_south_data -> terminal_south_0:data
	wire         node_131072_output_south_ready;         // terminal_south_0:ready -> node_131072:output_south_ready
	wire         node_131072_output_south_startofpacket; // node_131072:output_south_startofpacket -> terminal_south_0:startofpacket
	wire         node_131072_output_south_endofpacket;   // node_131072:output_south_endofpacket -> terminal_south_0:endofpacket
	wire   [1:0] node_131072_output_south_empty;         // node_131072:output_south_empty -> terminal_south_0:empty
	wire         node_131073_output_south_valid;         // node_131073:output_south_valid -> terminal_south_1:valid
	wire  [31:0] node_131073_output_south_data;          // node_131073:output_south_data -> terminal_south_1:data
	wire         node_131073_output_south_ready;         // terminal_south_1:ready -> node_131073:output_south_ready
	wire         node_131073_output_south_startofpacket; // node_131073:output_south_startofpacket -> terminal_south_1:startofpacket
	wire         node_131073_output_south_endofpacket;   // node_131073:output_south_endofpacket -> terminal_south_1:endofpacket
	wire   [1:0] node_131073_output_south_empty;         // node_131073:output_south_empty -> terminal_south_1:empty
	wire         node_131074_output_south_valid;         // node_131074:output_south_valid -> terminal_south_2:valid
	wire  [31:0] node_131074_output_south_data;          // node_131074:output_south_data -> terminal_south_2:data
	wire         node_131074_output_south_ready;         // terminal_south_2:ready -> node_131074:output_south_ready
	wire         node_131074_output_south_startofpacket; // node_131074:output_south_startofpacket -> terminal_south_2:startofpacket
	wire         node_131074_output_south_endofpacket;   // node_131074:output_south_endofpacket -> terminal_south_2:endofpacket
	wire   [1:0] node_131074_output_south_empty;         // node_131074:output_south_empty -> terminal_south_2:empty
	wire         node_131080_output_south_valid;         // node_131080:output_south_valid -> terminal_south_8:valid
	wire  [31:0] node_131080_output_south_data;          // node_131080:output_south_data -> terminal_south_8:data
	wire         node_131080_output_south_ready;         // terminal_south_8:ready -> node_131080:output_south_ready
	wire         node_131080_output_south_startofpacket; // node_131080:output_south_startofpacket -> terminal_south_8:startofpacket
	wire         node_131080_output_south_endofpacket;   // node_131080:output_south_endofpacket -> terminal_south_8:endofpacket
	wire   [1:0] node_131080_output_south_empty;         // node_131080:output_south_empty -> terminal_south_8:empty
	wire         node_131079_output_south_valid;         // node_131079:output_south_valid -> terminal_south_7:valid
	wire  [31:0] node_131079_output_south_data;          // node_131079:output_south_data -> terminal_south_7:data
	wire         node_131079_output_south_ready;         // terminal_south_7:ready -> node_131079:output_south_ready
	wire         node_131079_output_south_startofpacket; // node_131079:output_south_startofpacket -> terminal_south_7:startofpacket
	wire         node_131079_output_south_endofpacket;   // node_131079:output_south_endofpacket -> terminal_south_7:endofpacket
	wire   [1:0] node_131079_output_south_empty;         // node_131079:output_south_empty -> terminal_south_7:empty
	wire         node_131078_output_south_valid;         // node_131078:output_south_valid -> terminal_south_6:valid
	wire  [31:0] node_131078_output_south_data;          // node_131078:output_south_data -> terminal_south_6:data
	wire         node_131078_output_south_ready;         // terminal_south_6:ready -> node_131078:output_south_ready
	wire         node_131078_output_south_startofpacket; // node_131078:output_south_startofpacket -> terminal_south_6:startofpacket
	wire         node_131078_output_south_endofpacket;   // node_131078:output_south_endofpacket -> terminal_south_6:endofpacket
	wire   [1:0] node_131078_output_south_empty;         // node_131078:output_south_empty -> terminal_south_6:empty
	wire         node_131077_output_south_valid;         // node_131077:output_south_valid -> terminal_south_5:valid
	wire  [31:0] node_131077_output_south_data;          // node_131077:output_south_data -> terminal_south_5:data
	wire         node_131077_output_south_ready;         // terminal_south_5:ready -> node_131077:output_south_ready
	wire         node_131077_output_south_startofpacket; // node_131077:output_south_startofpacket -> terminal_south_5:startofpacket
	wire         node_131077_output_south_endofpacket;   // node_131077:output_south_endofpacket -> terminal_south_5:endofpacket
	wire   [1:0] node_131077_output_south_empty;         // node_131077:output_south_empty -> terminal_south_5:empty
	wire         node_131076_output_south_valid;         // node_131076:output_south_valid -> terminal_south_4:valid
	wire  [31:0] node_131076_output_south_data;          // node_131076:output_south_data -> terminal_south_4:data
	wire         node_131076_output_south_ready;         // terminal_south_4:ready -> node_131076:output_south_ready
	wire         node_131076_output_south_startofpacket; // node_131076:output_south_startofpacket -> terminal_south_4:startofpacket
	wire         node_131076_output_south_endofpacket;   // node_131076:output_south_endofpacket -> terminal_south_4:endofpacket
	wire   [1:0] node_131076_output_south_empty;         // node_131076:output_south_empty -> terminal_south_4:empty
	wire         node_131075_output_south_valid;         // node_131075:output_south_valid -> terminal_south_3:valid
	wire  [31:0] node_131075_output_south_data;          // node_131075:output_south_data -> terminal_south_3:data
	wire         node_131075_output_south_ready;         // terminal_south_3:ready -> node_131075:output_south_ready
	wire         node_131075_output_south_startofpacket; // node_131075:output_south_startofpacket -> terminal_south_3:startofpacket
	wire         node_131075_output_south_endofpacket;   // node_131075:output_south_endofpacket -> terminal_south_3:endofpacket
	wire   [1:0] node_131075_output_south_empty;         // node_131075:output_south_empty -> terminal_south_3:empty
	wire         node_1_output_west_valid;               // node_1:output_west_valid -> node_0:input_east_valid
	wire  [31:0] node_1_output_west_data;                // node_1:output_west_data -> node_0:input_east_data
	wire         node_1_output_west_ready;               // node_0:input_east_ready -> node_1:output_west_ready
	wire         node_1_output_west_startofpacket;       // node_1:output_west_startofpacket -> node_0:input_east_startofpacket
	wire         node_1_output_west_endofpacket;         // node_1:output_west_endofpacket -> node_0:input_east_endofpacket
	wire   [1:0] node_1_output_west_empty;               // node_1:output_west_empty -> node_0:input_east_empty
	wire         node_2_output_west_valid;               // node_2:output_west_valid -> node_1:input_east_valid
	wire  [31:0] node_2_output_west_data;                // node_2:output_west_data -> node_1:input_east_data
	wire         node_2_output_west_ready;               // node_1:input_east_ready -> node_2:output_west_ready
	wire         node_2_output_west_startofpacket;       // node_2:output_west_startofpacket -> node_1:input_east_startofpacket
	wire         node_2_output_west_endofpacket;         // node_2:output_west_endofpacket -> node_1:input_east_endofpacket
	wire   [1:0] node_2_output_west_empty;               // node_2:output_west_empty -> node_1:input_east_empty
	wire         node_65537_output_west_valid;           // node_65537:output_west_valid -> node_65536:input_east_valid
	wire  [31:0] node_65537_output_west_data;            // node_65537:output_west_data -> node_65536:input_east_data
	wire         node_65537_output_west_ready;           // node_65536:input_east_ready -> node_65537:output_west_ready
	wire         node_65537_output_west_startofpacket;   // node_65537:output_west_startofpacket -> node_65536:input_east_startofpacket
	wire         node_65537_output_west_endofpacket;     // node_65537:output_west_endofpacket -> node_65536:input_east_endofpacket
	wire   [1:0] node_65537_output_west_empty;           // node_65537:output_west_empty -> node_65536:input_east_empty
	wire         node_65538_output_west_valid;           // node_65538:output_west_valid -> node_65537:input_east_valid
	wire  [31:0] node_65538_output_west_data;            // node_65538:output_west_data -> node_65537:input_east_data
	wire         node_65538_output_west_ready;           // node_65537:input_east_ready -> node_65538:output_west_ready
	wire         node_65538_output_west_startofpacket;   // node_65538:output_west_startofpacket -> node_65537:input_east_startofpacket
	wire         node_65538_output_west_endofpacket;     // node_65538:output_west_endofpacket -> node_65537:input_east_endofpacket
	wire   [1:0] node_65538_output_west_empty;           // node_65538:output_west_empty -> node_65537:input_east_empty
	wire         node_131073_output_west_valid;          // node_131073:output_west_valid -> node_131072:input_east_valid
	wire  [31:0] node_131073_output_west_data;           // node_131073:output_west_data -> node_131072:input_east_data
	wire         node_131073_output_west_ready;          // node_131072:input_east_ready -> node_131073:output_west_ready
	wire         node_131073_output_west_startofpacket;  // node_131073:output_west_startofpacket -> node_131072:input_east_startofpacket
	wire         node_131073_output_west_endofpacket;    // node_131073:output_west_endofpacket -> node_131072:input_east_endofpacket
	wire   [1:0] node_131073_output_west_empty;          // node_131073:output_west_empty -> node_131072:input_east_empty
	wire         node_131074_output_west_valid;          // node_131074:output_west_valid -> node_131073:input_east_valid
	wire  [31:0] node_131074_output_west_data;           // node_131074:output_west_data -> node_131073:input_east_data
	wire         node_131074_output_west_ready;          // node_131073:input_east_ready -> node_131074:output_west_ready
	wire         node_131074_output_west_startofpacket;  // node_131074:output_west_startofpacket -> node_131073:input_east_startofpacket
	wire         node_131074_output_west_endofpacket;    // node_131074:output_west_endofpacket -> node_131073:input_east_endofpacket
	wire   [1:0] node_131074_output_west_empty;          // node_131074:output_west_empty -> node_131073:input_east_empty
	wire         node_8_output_west_valid;               // node_8:output_west_valid -> node_7:input_east_valid
	wire  [31:0] node_8_output_west_data;                // node_8:output_west_data -> node_7:input_east_data
	wire         node_8_output_west_ready;               // node_7:input_east_ready -> node_8:output_west_ready
	wire         node_8_output_west_startofpacket;       // node_8:output_west_startofpacket -> node_7:input_east_startofpacket
	wire         node_8_output_west_endofpacket;         // node_8:output_west_endofpacket -> node_7:input_east_endofpacket
	wire   [1:0] node_8_output_west_empty;               // node_8:output_west_empty -> node_7:input_east_empty
	wire         node_7_output_west_valid;               // node_7:output_west_valid -> node_6:input_east_valid
	wire  [31:0] node_7_output_west_data;                // node_7:output_west_data -> node_6:input_east_data
	wire         node_7_output_west_ready;               // node_6:input_east_ready -> node_7:output_west_ready
	wire         node_7_output_west_startofpacket;       // node_7:output_west_startofpacket -> node_6:input_east_startofpacket
	wire         node_7_output_west_endofpacket;         // node_7:output_west_endofpacket -> node_6:input_east_endofpacket
	wire   [1:0] node_7_output_west_empty;               // node_7:output_west_empty -> node_6:input_east_empty
	wire         node_6_output_west_valid;               // node_6:output_west_valid -> node_5:input_east_valid
	wire  [31:0] node_6_output_west_data;                // node_6:output_west_data -> node_5:input_east_data
	wire         node_6_output_west_ready;               // node_5:input_east_ready -> node_6:output_west_ready
	wire         node_6_output_west_startofpacket;       // node_6:output_west_startofpacket -> node_5:input_east_startofpacket
	wire         node_6_output_west_endofpacket;         // node_6:output_west_endofpacket -> node_5:input_east_endofpacket
	wire   [1:0] node_6_output_west_empty;               // node_6:output_west_empty -> node_5:input_east_empty
	wire         node_5_output_west_valid;               // node_5:output_west_valid -> node_4:input_east_valid
	wire  [31:0] node_5_output_west_data;                // node_5:output_west_data -> node_4:input_east_data
	wire         node_5_output_west_ready;               // node_4:input_east_ready -> node_5:output_west_ready
	wire         node_5_output_west_startofpacket;       // node_5:output_west_startofpacket -> node_4:input_east_startofpacket
	wire         node_5_output_west_endofpacket;         // node_5:output_west_endofpacket -> node_4:input_east_endofpacket
	wire   [1:0] node_5_output_west_empty;               // node_5:output_west_empty -> node_4:input_east_empty
	wire         node_4_output_west_valid;               // node_4:output_west_valid -> node_3:input_east_valid
	wire  [31:0] node_4_output_west_data;                // node_4:output_west_data -> node_3:input_east_data
	wire         node_4_output_west_ready;               // node_3:input_east_ready -> node_4:output_west_ready
	wire         node_4_output_west_startofpacket;       // node_4:output_west_startofpacket -> node_3:input_east_startofpacket
	wire         node_4_output_west_endofpacket;         // node_4:output_west_endofpacket -> node_3:input_east_endofpacket
	wire   [1:0] node_4_output_west_empty;               // node_4:output_west_empty -> node_3:input_east_empty
	wire         node_3_output_west_valid;               // node_3:output_west_valid -> node_2:input_east_valid
	wire  [31:0] node_3_output_west_data;                // node_3:output_west_data -> node_2:input_east_data
	wire         node_3_output_west_ready;               // node_2:input_east_ready -> node_3:output_west_ready
	wire         node_3_output_west_startofpacket;       // node_3:output_west_startofpacket -> node_2:input_east_startofpacket
	wire         node_3_output_west_endofpacket;         // node_3:output_west_endofpacket -> node_2:input_east_endofpacket
	wire   [1:0] node_3_output_west_empty;               // node_3:output_west_empty -> node_2:input_east_empty
	wire         node_65544_output_west_valid;           // node_65544:output_west_valid -> node_65543:input_east_valid
	wire  [31:0] node_65544_output_west_data;            // node_65544:output_west_data -> node_65543:input_east_data
	wire         node_65544_output_west_ready;           // node_65543:input_east_ready -> node_65544:output_west_ready
	wire         node_65544_output_west_startofpacket;   // node_65544:output_west_startofpacket -> node_65543:input_east_startofpacket
	wire         node_65544_output_west_endofpacket;     // node_65544:output_west_endofpacket -> node_65543:input_east_endofpacket
	wire   [1:0] node_65544_output_west_empty;           // node_65544:output_west_empty -> node_65543:input_east_empty
	wire         node_65543_output_west_valid;           // node_65543:output_west_valid -> node_65542:input_east_valid
	wire  [31:0] node_65543_output_west_data;            // node_65543:output_west_data -> node_65542:input_east_data
	wire         node_65543_output_west_ready;           // node_65542:input_east_ready -> node_65543:output_west_ready
	wire         node_65543_output_west_startofpacket;   // node_65543:output_west_startofpacket -> node_65542:input_east_startofpacket
	wire         node_65543_output_west_endofpacket;     // node_65543:output_west_endofpacket -> node_65542:input_east_endofpacket
	wire   [1:0] node_65543_output_west_empty;           // node_65543:output_west_empty -> node_65542:input_east_empty
	wire         node_65542_output_west_valid;           // node_65542:output_west_valid -> node_65541:input_east_valid
	wire  [31:0] node_65542_output_west_data;            // node_65542:output_west_data -> node_65541:input_east_data
	wire         node_65542_output_west_ready;           // node_65541:input_east_ready -> node_65542:output_west_ready
	wire         node_65542_output_west_startofpacket;   // node_65542:output_west_startofpacket -> node_65541:input_east_startofpacket
	wire         node_65542_output_west_endofpacket;     // node_65542:output_west_endofpacket -> node_65541:input_east_endofpacket
	wire   [1:0] node_65542_output_west_empty;           // node_65542:output_west_empty -> node_65541:input_east_empty
	wire         node_65541_output_west_valid;           // node_65541:output_west_valid -> node_65540:input_east_valid
	wire  [31:0] node_65541_output_west_data;            // node_65541:output_west_data -> node_65540:input_east_data
	wire         node_65541_output_west_ready;           // node_65540:input_east_ready -> node_65541:output_west_ready
	wire         node_65541_output_west_startofpacket;   // node_65541:output_west_startofpacket -> node_65540:input_east_startofpacket
	wire         node_65541_output_west_endofpacket;     // node_65541:output_west_endofpacket -> node_65540:input_east_endofpacket
	wire   [1:0] node_65541_output_west_empty;           // node_65541:output_west_empty -> node_65540:input_east_empty
	wire         node_65540_output_west_valid;           // node_65540:output_west_valid -> node_65539:input_east_valid
	wire  [31:0] node_65540_output_west_data;            // node_65540:output_west_data -> node_65539:input_east_data
	wire         node_65540_output_west_ready;           // node_65539:input_east_ready -> node_65540:output_west_ready
	wire         node_65540_output_west_startofpacket;   // node_65540:output_west_startofpacket -> node_65539:input_east_startofpacket
	wire         node_65540_output_west_endofpacket;     // node_65540:output_west_endofpacket -> node_65539:input_east_endofpacket
	wire   [1:0] node_65540_output_west_empty;           // node_65540:output_west_empty -> node_65539:input_east_empty
	wire         node_65539_output_west_valid;           // node_65539:output_west_valid -> node_65538:input_east_valid
	wire  [31:0] node_65539_output_west_data;            // node_65539:output_west_data -> node_65538:input_east_data
	wire         node_65539_output_west_ready;           // node_65538:input_east_ready -> node_65539:output_west_ready
	wire         node_65539_output_west_startofpacket;   // node_65539:output_west_startofpacket -> node_65538:input_east_startofpacket
	wire         node_65539_output_west_endofpacket;     // node_65539:output_west_endofpacket -> node_65538:input_east_endofpacket
	wire   [1:0] node_65539_output_west_empty;           // node_65539:output_west_empty -> node_65538:input_east_empty
	wire         node_131080_output_west_valid;          // node_131080:output_west_valid -> node_131079:input_east_valid
	wire  [31:0] node_131080_output_west_data;           // node_131080:output_west_data -> node_131079:input_east_data
	wire         node_131080_output_west_ready;          // node_131079:input_east_ready -> node_131080:output_west_ready
	wire         node_131080_output_west_startofpacket;  // node_131080:output_west_startofpacket -> node_131079:input_east_startofpacket
	wire         node_131080_output_west_endofpacket;    // node_131080:output_west_endofpacket -> node_131079:input_east_endofpacket
	wire   [1:0] node_131080_output_west_empty;          // node_131080:output_west_empty -> node_131079:input_east_empty
	wire         node_131079_output_west_valid;          // node_131079:output_west_valid -> node_131078:input_east_valid
	wire  [31:0] node_131079_output_west_data;           // node_131079:output_west_data -> node_131078:input_east_data
	wire         node_131079_output_west_ready;          // node_131078:input_east_ready -> node_131079:output_west_ready
	wire         node_131079_output_west_startofpacket;  // node_131079:output_west_startofpacket -> node_131078:input_east_startofpacket
	wire         node_131079_output_west_endofpacket;    // node_131079:output_west_endofpacket -> node_131078:input_east_endofpacket
	wire   [1:0] node_131079_output_west_empty;          // node_131079:output_west_empty -> node_131078:input_east_empty
	wire         node_131078_output_west_valid;          // node_131078:output_west_valid -> node_131077:input_east_valid
	wire  [31:0] node_131078_output_west_data;           // node_131078:output_west_data -> node_131077:input_east_data
	wire         node_131078_output_west_ready;          // node_131077:input_east_ready -> node_131078:output_west_ready
	wire         node_131078_output_west_startofpacket;  // node_131078:output_west_startofpacket -> node_131077:input_east_startofpacket
	wire         node_131078_output_west_endofpacket;    // node_131078:output_west_endofpacket -> node_131077:input_east_endofpacket
	wire   [1:0] node_131078_output_west_empty;          // node_131078:output_west_empty -> node_131077:input_east_empty
	wire         node_131077_output_west_valid;          // node_131077:output_west_valid -> node_131076:input_east_valid
	wire  [31:0] node_131077_output_west_data;           // node_131077:output_west_data -> node_131076:input_east_data
	wire         node_131077_output_west_ready;          // node_131076:input_east_ready -> node_131077:output_west_ready
	wire         node_131077_output_west_startofpacket;  // node_131077:output_west_startofpacket -> node_131076:input_east_startofpacket
	wire         node_131077_output_west_endofpacket;    // node_131077:output_west_endofpacket -> node_131076:input_east_endofpacket
	wire   [1:0] node_131077_output_west_empty;          // node_131077:output_west_empty -> node_131076:input_east_empty
	wire         node_131076_output_west_valid;          // node_131076:output_west_valid -> node_131075:input_east_valid
	wire  [31:0] node_131076_output_west_data;           // node_131076:output_west_data -> node_131075:input_east_data
	wire         node_131076_output_west_ready;          // node_131075:input_east_ready -> node_131076:output_west_ready
	wire         node_131076_output_west_startofpacket;  // node_131076:output_west_startofpacket -> node_131075:input_east_startofpacket
	wire         node_131076_output_west_endofpacket;    // node_131076:output_west_endofpacket -> node_131075:input_east_endofpacket
	wire   [1:0] node_131076_output_west_empty;          // node_131076:output_west_empty -> node_131075:input_east_empty
	wire         node_131075_output_west_valid;          // node_131075:output_west_valid -> node_131074:input_east_valid
	wire  [31:0] node_131075_output_west_data;           // node_131075:output_west_data -> node_131074:input_east_data
	wire         node_131075_output_west_ready;          // node_131074:input_east_ready -> node_131075:output_west_ready
	wire         node_131075_output_west_startofpacket;  // node_131075:output_west_startofpacket -> node_131074:input_east_startofpacket
	wire         node_131075_output_west_endofpacket;    // node_131075:output_west_endofpacket -> node_131074:input_east_endofpacket
	wire   [1:0] node_131075_output_west_empty;          // node_131075:output_west_empty -> node_131074:input_east_empty
	wire         node_0_output_west_valid;               // node_0:output_west_valid -> terminal_west_0:valid
	wire  [31:0] node_0_output_west_data;                // node_0:output_west_data -> terminal_west_0:data
	wire         node_0_output_west_ready;               // terminal_west_0:ready -> node_0:output_west_ready
	wire         node_0_output_west_startofpacket;       // node_0:output_west_startofpacket -> terminal_west_0:startofpacket
	wire         node_0_output_west_endofpacket;         // node_0:output_west_endofpacket -> terminal_west_0:endofpacket
	wire   [1:0] node_0_output_west_empty;               // node_0:output_west_empty -> terminal_west_0:empty
	wire         node_65536_output_west_valid;           // node_65536:output_west_valid -> terminal_west_1:valid
	wire  [31:0] node_65536_output_west_data;            // node_65536:output_west_data -> terminal_west_1:data
	wire         node_65536_output_west_ready;           // terminal_west_1:ready -> node_65536:output_west_ready
	wire         node_65536_output_west_startofpacket;   // node_65536:output_west_startofpacket -> terminal_west_1:startofpacket
	wire         node_65536_output_west_endofpacket;     // node_65536:output_west_endofpacket -> terminal_west_1:endofpacket
	wire   [1:0] node_65536_output_west_empty;           // node_65536:output_west_empty -> terminal_west_1:empty
	wire         node_131072_output_west_valid;          // node_131072:output_west_valid -> terminal_west_2:valid
	wire  [31:0] node_131072_output_west_data;           // node_131072:output_west_data -> terminal_west_2:data
	wire         node_131072_output_west_ready;          // terminal_west_2:ready -> node_131072:output_west_ready
	wire         node_131072_output_west_startofpacket;  // node_131072:output_west_startofpacket -> terminal_west_2:startofpacket
	wire         node_131072_output_west_endofpacket;    // node_131072:output_west_endofpacket -> terminal_west_2:endofpacket
	wire   [1:0] node_131072_output_west_empty;          // node_131072:output_west_empty -> terminal_west_2:empty
	wire         rst_controller_reset_out_reset;         // rst_controller:reset_out -> [terminal_east_0:reset_n, terminal_east_1:reset_n, terminal_east_2:reset_n, terminal_north_0:reset_n, terminal_north_1:reset_n, terminal_north_2:reset_n, terminal_north_3:reset_n, terminal_north_4:reset_n, terminal_north_5:reset_n, terminal_north_6:reset_n, terminal_north_7:reset_n, terminal_north_8:reset_n, terminal_south_0:reset_n, terminal_south_1:reset_n, terminal_south_2:reset_n, terminal_south_3:reset_n, terminal_south_4:reset_n, terminal_south_5:reset_n, terminal_south_6:reset_n, terminal_south_7:reset_n, terminal_south_8:reset_n, terminal_west_0:reset_n, terminal_west_1:reset_n, terminal_west_2:reset_n]

	dircc_system_rtl_gals_test_version_node_0 node_0 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_1_output_west_data),               //   input_east.data
		.input_east_valid           (node_1_output_west_valid),              //             .valid
		.input_east_ready           (node_1_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_1_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_1_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_1_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65536_output_north_data),          //  input_south.data
		.input_south_valid          (node_65536_output_north_valid),         //             .valid
		.input_south_ready          (node_65536_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65536_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65536_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65536_output_north_empty),         //             .empty
		.input_west_data            (),                                      //   input_west.data
		.input_west_valid           (),                                      //             .valid
		.input_west_ready           (),                                      //             .ready
		.input_west_startofpacket   (),                                      //             .startofpacket
		.input_west_endofpacket     (),                                      //             .endofpacket
		.input_west_empty           (),                                      //             .empty
		.mem_address                (node_0_mem_address),                    //          mem.address
		.mem_readdata               (node_0_mem_readdata),                   //             .readdata
		.mem_write                  (node_0_mem_write),                      //             .write
		.mem_writedata              (node_0_mem_writedata),                  //             .writedata
		.output_east_data           (node_0_output_east_data),               //  output_east.data
		.output_east_valid          (node_0_output_east_valid),              //             .valid
		.output_east_ready          (node_0_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_0_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_0_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_0_output_east_empty),              //             .empty
		.output_north_data          (node_0_output_north_data),              // output_north.data
		.output_north_valid         (node_0_output_north_valid),             //             .valid
		.output_north_ready         (node_0_output_north_ready),             //             .ready
		.output_north_startofpacket (node_0_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_0_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_0_output_north_empty),             //             .empty
		.output_south_data          (node_0_output_south_data),              // output_south.data
		.output_south_valid         (node_0_output_south_valid),             //             .valid
		.output_south_ready         (node_0_output_south_ready),             //             .ready
		.output_south_startofpacket (node_0_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_0_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_0_output_south_empty),             //             .empty
		.output_west_data           (node_0_output_west_data),               //  output_west.data
		.output_west_valid          (node_0_output_west_valid),              //             .valid
		.output_west_ready          (node_0_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_0_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_0_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_0_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_1 node_1 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_2_output_west_data),               //   input_east.data
		.input_east_valid           (node_2_output_west_valid),              //             .valid
		.input_east_ready           (node_2_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_2_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_2_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_2_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65537_output_north_data),          //  input_south.data
		.input_south_valid          (node_65537_output_north_valid),         //             .valid
		.input_south_ready          (node_65537_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65537_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65537_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65537_output_north_empty),         //             .empty
		.input_west_data            (node_0_output_east_data),               //   input_west.data
		.input_west_valid           (node_0_output_east_valid),              //             .valid
		.input_west_ready           (node_0_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_0_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_0_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_0_output_east_empty),              //             .empty
		.mem_address                (node_1_mem_address),                    //          mem.address
		.mem_readdata               (node_1_mem_readdata),                   //             .readdata
		.mem_write                  (node_1_mem_write),                      //             .write
		.mem_writedata              (node_1_mem_writedata),                  //             .writedata
		.output_east_data           (node_1_output_east_data),               //  output_east.data
		.output_east_valid          (node_1_output_east_valid),              //             .valid
		.output_east_ready          (node_1_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_1_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_1_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_1_output_east_empty),              //             .empty
		.output_north_data          (node_1_output_north_data),              // output_north.data
		.output_north_valid         (node_1_output_north_valid),             //             .valid
		.output_north_ready         (node_1_output_north_ready),             //             .ready
		.output_north_startofpacket (node_1_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_1_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_1_output_north_empty),             //             .empty
		.output_south_data          (node_1_output_south_data),              // output_south.data
		.output_south_valid         (node_1_output_south_valid),             //             .valid
		.output_south_ready         (node_1_output_south_ready),             //             .ready
		.output_south_startofpacket (node_1_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_1_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_1_output_south_empty),             //             .empty
		.output_west_data           (node_1_output_west_data),               //  output_west.data
		.output_west_valid          (node_1_output_west_valid),              //             .valid
		.output_west_ready          (node_1_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_1_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_1_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_1_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131072 node_131072 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131073_output_west_data),           //   input_east.data
		.input_east_valid           (node_131073_output_west_valid),          //             .valid
		.input_east_ready           (node_131073_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131073_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131073_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131073_output_west_empty),          //             .empty
		.input_north_data           (node_65536_output_south_data),           //  input_north.data
		.input_north_valid          (node_65536_output_south_valid),          //             .valid
		.input_north_ready          (node_65536_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65536_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65536_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65536_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (),                                       //   input_west.data
		.input_west_valid           (),                                       //             .valid
		.input_west_ready           (),                                       //             .ready
		.input_west_startofpacket   (),                                       //             .startofpacket
		.input_west_endofpacket     (),                                       //             .endofpacket
		.input_west_empty           (),                                       //             .empty
		.mem_address                (node_131072_mem_address),                //          mem.address
		.mem_readdata               (node_131072_mem_readdata),               //             .readdata
		.mem_write                  (node_131072_mem_write),                  //             .write
		.mem_writedata              (node_131072_mem_writedata),              //             .writedata
		.output_east_data           (node_131072_output_east_data),           //  output_east.data
		.output_east_valid          (node_131072_output_east_valid),          //             .valid
		.output_east_ready          (node_131072_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131072_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131072_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131072_output_east_empty),          //             .empty
		.output_north_data          (node_131072_output_north_data),          // output_north.data
		.output_north_valid         (node_131072_output_north_valid),         //             .valid
		.output_north_ready         (node_131072_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131072_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131072_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131072_output_north_empty),         //             .empty
		.output_south_data          (node_131072_output_south_data),          // output_south.data
		.output_south_valid         (node_131072_output_south_valid),         //             .valid
		.output_south_ready         (node_131072_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131072_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131072_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131072_output_south_empty),         //             .empty
		.output_west_data           (node_131072_output_west_data),           //  output_west.data
		.output_west_valid          (node_131072_output_west_valid),          //             .valid
		.output_west_ready          (node_131072_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131072_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131072_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131072_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131073 node_131073 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131074_output_west_data),           //   input_east.data
		.input_east_valid           (node_131074_output_west_valid),          //             .valid
		.input_east_ready           (node_131074_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131074_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131074_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131074_output_west_empty),          //             .empty
		.input_north_data           (node_65537_output_south_data),           //  input_north.data
		.input_north_valid          (node_65537_output_south_valid),          //             .valid
		.input_north_ready          (node_65537_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65537_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65537_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65537_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131072_output_east_data),           //   input_west.data
		.input_west_valid           (node_131072_output_east_valid),          //             .valid
		.input_west_ready           (node_131072_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131072_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131072_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131072_output_east_empty),          //             .empty
		.mem_address                (node_131073_mem_address),                //          mem.address
		.mem_readdata               (node_131073_mem_readdata),               //             .readdata
		.mem_write                  (node_131073_mem_write),                  //             .write
		.mem_writedata              (node_131073_mem_writedata),              //             .writedata
		.output_east_data           (node_131073_output_east_data),           //  output_east.data
		.output_east_valid          (node_131073_output_east_valid),          //             .valid
		.output_east_ready          (node_131073_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131073_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131073_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131073_output_east_empty),          //             .empty
		.output_north_data          (node_131073_output_north_data),          // output_north.data
		.output_north_valid         (node_131073_output_north_valid),         //             .valid
		.output_north_ready         (node_131073_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131073_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131073_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131073_output_north_empty),         //             .empty
		.output_south_data          (node_131073_output_south_data),          // output_south.data
		.output_south_valid         (node_131073_output_south_valid),         //             .valid
		.output_south_ready         (node_131073_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131073_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131073_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131073_output_south_empty),         //             .empty
		.output_west_data           (node_131073_output_west_data),           //  output_west.data
		.output_west_valid          (node_131073_output_west_valid),          //             .valid
		.output_west_ready          (node_131073_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131073_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131073_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131073_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131074 node_131074 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131075_output_west_data),           //   input_east.data
		.input_east_valid           (node_131075_output_west_valid),          //             .valid
		.input_east_ready           (node_131075_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131075_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131075_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131075_output_west_empty),          //             .empty
		.input_north_data           (node_65538_output_south_data),           //  input_north.data
		.input_north_valid          (node_65538_output_south_valid),          //             .valid
		.input_north_ready          (node_65538_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65538_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65538_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65538_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131073_output_east_data),           //   input_west.data
		.input_west_valid           (node_131073_output_east_valid),          //             .valid
		.input_west_ready           (node_131073_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131073_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131073_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131073_output_east_empty),          //             .empty
		.mem_address                (node_131074_mem_address),                //          mem.address
		.mem_readdata               (node_131074_mem_readdata),               //             .readdata
		.mem_write                  (node_131074_mem_write),                  //             .write
		.mem_writedata              (node_131074_mem_writedata),              //             .writedata
		.output_east_data           (node_131074_output_east_data),           //  output_east.data
		.output_east_valid          (node_131074_output_east_valid),          //             .valid
		.output_east_ready          (node_131074_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131074_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131074_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131074_output_east_empty),          //             .empty
		.output_north_data          (node_131074_output_north_data),          // output_north.data
		.output_north_valid         (node_131074_output_north_valid),         //             .valid
		.output_north_ready         (node_131074_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131074_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131074_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131074_output_north_empty),         //             .empty
		.output_south_data          (node_131074_output_south_data),          // output_south.data
		.output_south_valid         (node_131074_output_south_valid),         //             .valid
		.output_south_ready         (node_131074_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131074_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131074_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131074_output_south_empty),         //             .empty
		.output_west_data           (node_131074_output_west_data),           //  output_west.data
		.output_west_valid          (node_131074_output_west_valid),          //             .valid
		.output_west_ready          (node_131074_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131074_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131074_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131074_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131075 node_131075 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131076_output_west_data),           //   input_east.data
		.input_east_valid           (node_131076_output_west_valid),          //             .valid
		.input_east_ready           (node_131076_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131076_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131076_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131076_output_west_empty),          //             .empty
		.input_north_data           (node_65539_output_south_data),           //  input_north.data
		.input_north_valid          (node_65539_output_south_valid),          //             .valid
		.input_north_ready          (node_65539_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65539_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65539_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65539_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131074_output_east_data),           //   input_west.data
		.input_west_valid           (node_131074_output_east_valid),          //             .valid
		.input_west_ready           (node_131074_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131074_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131074_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131074_output_east_empty),          //             .empty
		.mem_address                (node_131075_mem_address),                //          mem.address
		.mem_readdata               (node_131075_mem_readdata),               //             .readdata
		.mem_write                  (node_131075_mem_write),                  //             .write
		.mem_writedata              (node_131075_mem_writedata),              //             .writedata
		.output_east_data           (node_131075_output_east_data),           //  output_east.data
		.output_east_valid          (node_131075_output_east_valid),          //             .valid
		.output_east_ready          (node_131075_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131075_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131075_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131075_output_east_empty),          //             .empty
		.output_north_data          (node_131075_output_north_data),          // output_north.data
		.output_north_valid         (node_131075_output_north_valid),         //             .valid
		.output_north_ready         (node_131075_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131075_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131075_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131075_output_north_empty),         //             .empty
		.output_south_data          (node_131075_output_south_data),          // output_south.data
		.output_south_valid         (node_131075_output_south_valid),         //             .valid
		.output_south_ready         (node_131075_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131075_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131075_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131075_output_south_empty),         //             .empty
		.output_west_data           (node_131075_output_west_data),           //  output_west.data
		.output_west_valid          (node_131075_output_west_valid),          //             .valid
		.output_west_ready          (node_131075_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131075_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131075_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131075_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131076 node_131076 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131077_output_west_data),           //   input_east.data
		.input_east_valid           (node_131077_output_west_valid),          //             .valid
		.input_east_ready           (node_131077_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131077_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131077_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131077_output_west_empty),          //             .empty
		.input_north_data           (node_65540_output_south_data),           //  input_north.data
		.input_north_valid          (node_65540_output_south_valid),          //             .valid
		.input_north_ready          (node_65540_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65540_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65540_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65540_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131075_output_east_data),           //   input_west.data
		.input_west_valid           (node_131075_output_east_valid),          //             .valid
		.input_west_ready           (node_131075_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131075_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131075_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131075_output_east_empty),          //             .empty
		.mem_address                (node_131076_mem_address),                //          mem.address
		.mem_readdata               (node_131076_mem_readdata),               //             .readdata
		.mem_write                  (node_131076_mem_write),                  //             .write
		.mem_writedata              (node_131076_mem_writedata),              //             .writedata
		.output_east_data           (node_131076_output_east_data),           //  output_east.data
		.output_east_valid          (node_131076_output_east_valid),          //             .valid
		.output_east_ready          (node_131076_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131076_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131076_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131076_output_east_empty),          //             .empty
		.output_north_data          (node_131076_output_north_data),          // output_north.data
		.output_north_valid         (node_131076_output_north_valid),         //             .valid
		.output_north_ready         (node_131076_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131076_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131076_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131076_output_north_empty),         //             .empty
		.output_south_data          (node_131076_output_south_data),          // output_south.data
		.output_south_valid         (node_131076_output_south_valid),         //             .valid
		.output_south_ready         (node_131076_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131076_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131076_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131076_output_south_empty),         //             .empty
		.output_west_data           (node_131076_output_west_data),           //  output_west.data
		.output_west_valid          (node_131076_output_west_valid),          //             .valid
		.output_west_ready          (node_131076_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131076_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131076_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131076_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131077 node_131077 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131078_output_west_data),           //   input_east.data
		.input_east_valid           (node_131078_output_west_valid),          //             .valid
		.input_east_ready           (node_131078_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131078_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131078_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131078_output_west_empty),          //             .empty
		.input_north_data           (node_65541_output_south_data),           //  input_north.data
		.input_north_valid          (node_65541_output_south_valid),          //             .valid
		.input_north_ready          (node_65541_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65541_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65541_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65541_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131076_output_east_data),           //   input_west.data
		.input_west_valid           (node_131076_output_east_valid),          //             .valid
		.input_west_ready           (node_131076_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131076_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131076_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131076_output_east_empty),          //             .empty
		.mem_address                (node_131077_mem_address),                //          mem.address
		.mem_readdata               (node_131077_mem_readdata),               //             .readdata
		.mem_write                  (node_131077_mem_write),                  //             .write
		.mem_writedata              (node_131077_mem_writedata),              //             .writedata
		.output_east_data           (node_131077_output_east_data),           //  output_east.data
		.output_east_valid          (node_131077_output_east_valid),          //             .valid
		.output_east_ready          (node_131077_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131077_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131077_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131077_output_east_empty),          //             .empty
		.output_north_data          (node_131077_output_north_data),          // output_north.data
		.output_north_valid         (node_131077_output_north_valid),         //             .valid
		.output_north_ready         (node_131077_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131077_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131077_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131077_output_north_empty),         //             .empty
		.output_south_data          (node_131077_output_south_data),          // output_south.data
		.output_south_valid         (node_131077_output_south_valid),         //             .valid
		.output_south_ready         (node_131077_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131077_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131077_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131077_output_south_empty),         //             .empty
		.output_west_data           (node_131077_output_west_data),           //  output_west.data
		.output_west_valid          (node_131077_output_west_valid),          //             .valid
		.output_west_ready          (node_131077_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131077_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131077_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131077_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131078 node_131078 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131079_output_west_data),           //   input_east.data
		.input_east_valid           (node_131079_output_west_valid),          //             .valid
		.input_east_ready           (node_131079_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131079_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131079_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131079_output_west_empty),          //             .empty
		.input_north_data           (node_65542_output_south_data),           //  input_north.data
		.input_north_valid          (node_65542_output_south_valid),          //             .valid
		.input_north_ready          (node_65542_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65542_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65542_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65542_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131077_output_east_data),           //   input_west.data
		.input_west_valid           (node_131077_output_east_valid),          //             .valid
		.input_west_ready           (node_131077_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131077_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131077_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131077_output_east_empty),          //             .empty
		.mem_address                (node_131078_mem_address),                //          mem.address
		.mem_readdata               (node_131078_mem_readdata),               //             .readdata
		.mem_write                  (node_131078_mem_write),                  //             .write
		.mem_writedata              (node_131078_mem_writedata),              //             .writedata
		.output_east_data           (node_131078_output_east_data),           //  output_east.data
		.output_east_valid          (node_131078_output_east_valid),          //             .valid
		.output_east_ready          (node_131078_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131078_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131078_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131078_output_east_empty),          //             .empty
		.output_north_data          (node_131078_output_north_data),          // output_north.data
		.output_north_valid         (node_131078_output_north_valid),         //             .valid
		.output_north_ready         (node_131078_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131078_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131078_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131078_output_north_empty),         //             .empty
		.output_south_data          (node_131078_output_south_data),          // output_south.data
		.output_south_valid         (node_131078_output_south_valid),         //             .valid
		.output_south_ready         (node_131078_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131078_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131078_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131078_output_south_empty),         //             .empty
		.output_west_data           (node_131078_output_west_data),           //  output_west.data
		.output_west_valid          (node_131078_output_west_valid),          //             .valid
		.output_west_ready          (node_131078_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131078_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131078_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131078_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131079 node_131079 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_131080_output_west_data),           //   input_east.data
		.input_east_valid           (node_131080_output_west_valid),          //             .valid
		.input_east_ready           (node_131080_output_west_ready),          //             .ready
		.input_east_startofpacket   (node_131080_output_west_startofpacket),  //             .startofpacket
		.input_east_endofpacket     (node_131080_output_west_endofpacket),    //             .endofpacket
		.input_east_empty           (node_131080_output_west_empty),          //             .empty
		.input_north_data           (node_65543_output_south_data),           //  input_north.data
		.input_north_valid          (node_65543_output_south_valid),          //             .valid
		.input_north_ready          (node_65543_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65543_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65543_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65543_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131078_output_east_data),           //   input_west.data
		.input_west_valid           (node_131078_output_east_valid),          //             .valid
		.input_west_ready           (node_131078_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131078_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131078_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131078_output_east_empty),          //             .empty
		.mem_address                (node_131079_mem_address),                //          mem.address
		.mem_readdata               (node_131079_mem_readdata),               //             .readdata
		.mem_write                  (node_131079_mem_write),                  //             .write
		.mem_writedata              (node_131079_mem_writedata),              //             .writedata
		.output_east_data           (node_131079_output_east_data),           //  output_east.data
		.output_east_valid          (node_131079_output_east_valid),          //             .valid
		.output_east_ready          (node_131079_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131079_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131079_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131079_output_east_empty),          //             .empty
		.output_north_data          (node_131079_output_north_data),          // output_north.data
		.output_north_valid         (node_131079_output_north_valid),         //             .valid
		.output_north_ready         (node_131079_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131079_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131079_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131079_output_north_empty),         //             .empty
		.output_south_data          (node_131079_output_south_data),          // output_south.data
		.output_south_valid         (node_131079_output_south_valid),         //             .valid
		.output_south_ready         (node_131079_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131079_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131079_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131079_output_south_empty),         //             .empty
		.output_west_data           (node_131079_output_west_data),           //  output_west.data
		.output_west_valid          (node_131079_output_west_valid),          //             .valid
		.output_west_ready          (node_131079_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131079_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131079_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131079_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_131080 node_131080 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (),                                       //   input_east.data
		.input_east_valid           (),                                       //             .valid
		.input_east_ready           (),                                       //             .ready
		.input_east_startofpacket   (),                                       //             .startofpacket
		.input_east_endofpacket     (),                                       //             .endofpacket
		.input_east_empty           (),                                       //             .empty
		.input_north_data           (node_65544_output_south_data),           //  input_north.data
		.input_north_valid          (node_65544_output_south_valid),          //             .valid
		.input_north_ready          (node_65544_output_south_ready),          //             .ready
		.input_north_startofpacket  (node_65544_output_south_startofpacket),  //             .startofpacket
		.input_north_endofpacket    (node_65544_output_south_endofpacket),    //             .endofpacket
		.input_north_empty          (node_65544_output_south_empty),          //             .empty
		.input_south_data           (),                                       //  input_south.data
		.input_south_valid          (),                                       //             .valid
		.input_south_ready          (),                                       //             .ready
		.input_south_startofpacket  (),                                       //             .startofpacket
		.input_south_endofpacket    (),                                       //             .endofpacket
		.input_south_empty          (),                                       //             .empty
		.input_west_data            (node_131079_output_east_data),           //   input_west.data
		.input_west_valid           (node_131079_output_east_valid),          //             .valid
		.input_west_ready           (node_131079_output_east_ready),          //             .ready
		.input_west_startofpacket   (node_131079_output_east_startofpacket),  //             .startofpacket
		.input_west_endofpacket     (node_131079_output_east_endofpacket),    //             .endofpacket
		.input_west_empty           (node_131079_output_east_empty),          //             .empty
		.mem_address                (node_131080_mem_address),                //          mem.address
		.mem_readdata               (node_131080_mem_readdata),               //             .readdata
		.mem_write                  (node_131080_mem_write),                  //             .write
		.mem_writedata              (node_131080_mem_writedata),              //             .writedata
		.output_east_data           (node_131080_output_east_data),           //  output_east.data
		.output_east_valid          (node_131080_output_east_valid),          //             .valid
		.output_east_ready          (node_131080_output_east_ready),          //             .ready
		.output_east_startofpacket  (node_131080_output_east_startofpacket),  //             .startofpacket
		.output_east_endofpacket    (node_131080_output_east_endofpacket),    //             .endofpacket
		.output_east_empty          (node_131080_output_east_empty),          //             .empty
		.output_north_data          (node_131080_output_north_data),          // output_north.data
		.output_north_valid         (node_131080_output_north_valid),         //             .valid
		.output_north_ready         (node_131080_output_north_ready),         //             .ready
		.output_north_startofpacket (node_131080_output_north_startofpacket), //             .startofpacket
		.output_north_endofpacket   (node_131080_output_north_endofpacket),   //             .endofpacket
		.output_north_empty         (node_131080_output_north_empty),         //             .empty
		.output_south_data          (node_131080_output_south_data),          // output_south.data
		.output_south_valid         (node_131080_output_south_valid),         //             .valid
		.output_south_ready         (node_131080_output_south_ready),         //             .ready
		.output_south_startofpacket (node_131080_output_south_startofpacket), //             .startofpacket
		.output_south_endofpacket   (node_131080_output_south_endofpacket),   //             .endofpacket
		.output_south_empty         (node_131080_output_south_empty),         //             .empty
		.output_west_data           (node_131080_output_west_data),           //  output_west.data
		.output_west_valid          (node_131080_output_west_valid),          //             .valid
		.output_west_ready          (node_131080_output_west_ready),          //             .ready
		.output_west_startofpacket  (node_131080_output_west_startofpacket),  //             .startofpacket
		.output_west_endofpacket    (node_131080_output_west_endofpacket),    //             .endofpacket
		.output_west_empty          (node_131080_output_west_empty),          //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_2 node_2 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_3_output_west_data),               //   input_east.data
		.input_east_valid           (node_3_output_west_valid),              //             .valid
		.input_east_ready           (node_3_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_3_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_3_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_3_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65538_output_north_data),          //  input_south.data
		.input_south_valid          (node_65538_output_north_valid),         //             .valid
		.input_south_ready          (node_65538_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65538_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65538_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65538_output_north_empty),         //             .empty
		.input_west_data            (node_1_output_east_data),               //   input_west.data
		.input_west_valid           (node_1_output_east_valid),              //             .valid
		.input_west_ready           (node_1_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_1_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_1_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_1_output_east_empty),              //             .empty
		.mem_address                (node_2_mem_address),                    //          mem.address
		.mem_readdata               (node_2_mem_readdata),                   //             .readdata
		.mem_write                  (node_2_mem_write),                      //             .write
		.mem_writedata              (node_2_mem_writedata),                  //             .writedata
		.output_east_data           (node_2_output_east_data),               //  output_east.data
		.output_east_valid          (node_2_output_east_valid),              //             .valid
		.output_east_ready          (node_2_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_2_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_2_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_2_output_east_empty),              //             .empty
		.output_north_data          (node_2_output_north_data),              // output_north.data
		.output_north_valid         (node_2_output_north_valid),             //             .valid
		.output_north_ready         (node_2_output_north_ready),             //             .ready
		.output_north_startofpacket (node_2_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_2_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_2_output_north_empty),             //             .empty
		.output_south_data          (node_2_output_south_data),              // output_south.data
		.output_south_valid         (node_2_output_south_valid),             //             .valid
		.output_south_ready         (node_2_output_south_ready),             //             .ready
		.output_south_startofpacket (node_2_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_2_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_2_output_south_empty),             //             .empty
		.output_west_data           (node_2_output_west_data),               //  output_west.data
		.output_west_valid          (node_2_output_west_valid),              //             .valid
		.output_west_ready          (node_2_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_2_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_2_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_2_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_3 node_3 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_4_output_west_data),               //   input_east.data
		.input_east_valid           (node_4_output_west_valid),              //             .valid
		.input_east_ready           (node_4_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_4_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_4_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_4_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65539_output_north_data),          //  input_south.data
		.input_south_valid          (node_65539_output_north_valid),         //             .valid
		.input_south_ready          (node_65539_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65539_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65539_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65539_output_north_empty),         //             .empty
		.input_west_data            (node_2_output_east_data),               //   input_west.data
		.input_west_valid           (node_2_output_east_valid),              //             .valid
		.input_west_ready           (node_2_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_2_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_2_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_2_output_east_empty),              //             .empty
		.mem_address                (node_3_mem_address),                    //          mem.address
		.mem_readdata               (node_3_mem_readdata),                   //             .readdata
		.mem_write                  (node_3_mem_write),                      //             .write
		.mem_writedata              (node_3_mem_writedata),                  //             .writedata
		.output_east_data           (node_3_output_east_data),               //  output_east.data
		.output_east_valid          (node_3_output_east_valid),              //             .valid
		.output_east_ready          (node_3_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_3_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_3_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_3_output_east_empty),              //             .empty
		.output_north_data          (node_3_output_north_data),              // output_north.data
		.output_north_valid         (node_3_output_north_valid),             //             .valid
		.output_north_ready         (node_3_output_north_ready),             //             .ready
		.output_north_startofpacket (node_3_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_3_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_3_output_north_empty),             //             .empty
		.output_south_data          (node_3_output_south_data),              // output_south.data
		.output_south_valid         (node_3_output_south_valid),             //             .valid
		.output_south_ready         (node_3_output_south_ready),             //             .ready
		.output_south_startofpacket (node_3_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_3_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_3_output_south_empty),             //             .empty
		.output_west_data           (node_3_output_west_data),               //  output_west.data
		.output_west_valid          (node_3_output_west_valid),              //             .valid
		.output_west_ready          (node_3_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_3_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_3_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_3_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_4 node_4 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_5_output_west_data),               //   input_east.data
		.input_east_valid           (node_5_output_west_valid),              //             .valid
		.input_east_ready           (node_5_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_5_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_5_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_5_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65540_output_north_data),          //  input_south.data
		.input_south_valid          (node_65540_output_north_valid),         //             .valid
		.input_south_ready          (node_65540_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65540_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65540_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65540_output_north_empty),         //             .empty
		.input_west_data            (node_3_output_east_data),               //   input_west.data
		.input_west_valid           (node_3_output_east_valid),              //             .valid
		.input_west_ready           (node_3_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_3_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_3_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_3_output_east_empty),              //             .empty
		.mem_address                (node_4_mem_address),                    //          mem.address
		.mem_readdata               (node_4_mem_readdata),                   //             .readdata
		.mem_write                  (node_4_mem_write),                      //             .write
		.mem_writedata              (node_4_mem_writedata),                  //             .writedata
		.output_east_data           (node_4_output_east_data),               //  output_east.data
		.output_east_valid          (node_4_output_east_valid),              //             .valid
		.output_east_ready          (node_4_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_4_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_4_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_4_output_east_empty),              //             .empty
		.output_north_data          (node_4_output_north_data),              // output_north.data
		.output_north_valid         (node_4_output_north_valid),             //             .valid
		.output_north_ready         (node_4_output_north_ready),             //             .ready
		.output_north_startofpacket (node_4_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_4_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_4_output_north_empty),             //             .empty
		.output_south_data          (node_4_output_south_data),              // output_south.data
		.output_south_valid         (node_4_output_south_valid),             //             .valid
		.output_south_ready         (node_4_output_south_ready),             //             .ready
		.output_south_startofpacket (node_4_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_4_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_4_output_south_empty),             //             .empty
		.output_west_data           (node_4_output_west_data),               //  output_west.data
		.output_west_valid          (node_4_output_west_valid),              //             .valid
		.output_west_ready          (node_4_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_4_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_4_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_4_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_5 node_5 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_6_output_west_data),               //   input_east.data
		.input_east_valid           (node_6_output_west_valid),              //             .valid
		.input_east_ready           (node_6_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_6_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_6_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_6_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65541_output_north_data),          //  input_south.data
		.input_south_valid          (node_65541_output_north_valid),         //             .valid
		.input_south_ready          (node_65541_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65541_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65541_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65541_output_north_empty),         //             .empty
		.input_west_data            (node_4_output_east_data),               //   input_west.data
		.input_west_valid           (node_4_output_east_valid),              //             .valid
		.input_west_ready           (node_4_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_4_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_4_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_4_output_east_empty),              //             .empty
		.mem_address                (node_5_mem_address),                    //          mem.address
		.mem_readdata               (node_5_mem_readdata),                   //             .readdata
		.mem_write                  (node_5_mem_write),                      //             .write
		.mem_writedata              (node_5_mem_writedata),                  //             .writedata
		.output_east_data           (node_5_output_east_data),               //  output_east.data
		.output_east_valid          (node_5_output_east_valid),              //             .valid
		.output_east_ready          (node_5_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_5_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_5_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_5_output_east_empty),              //             .empty
		.output_north_data          (node_5_output_north_data),              // output_north.data
		.output_north_valid         (node_5_output_north_valid),             //             .valid
		.output_north_ready         (node_5_output_north_ready),             //             .ready
		.output_north_startofpacket (node_5_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_5_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_5_output_north_empty),             //             .empty
		.output_south_data          (node_5_output_south_data),              // output_south.data
		.output_south_valid         (node_5_output_south_valid),             //             .valid
		.output_south_ready         (node_5_output_south_ready),             //             .ready
		.output_south_startofpacket (node_5_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_5_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_5_output_south_empty),             //             .empty
		.output_west_data           (node_5_output_west_data),               //  output_west.data
		.output_west_valid          (node_5_output_west_valid),              //             .valid
		.output_west_ready          (node_5_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_5_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_5_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_5_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_6 node_6 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_7_output_west_data),               //   input_east.data
		.input_east_valid           (node_7_output_west_valid),              //             .valid
		.input_east_ready           (node_7_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_7_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_7_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_7_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65542_output_north_data),          //  input_south.data
		.input_south_valid          (node_65542_output_north_valid),         //             .valid
		.input_south_ready          (node_65542_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65542_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65542_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65542_output_north_empty),         //             .empty
		.input_west_data            (node_5_output_east_data),               //   input_west.data
		.input_west_valid           (node_5_output_east_valid),              //             .valid
		.input_west_ready           (node_5_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_5_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_5_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_5_output_east_empty),              //             .empty
		.mem_address                (node_6_mem_address),                    //          mem.address
		.mem_readdata               (node_6_mem_readdata),                   //             .readdata
		.mem_write                  (node_6_mem_write),                      //             .write
		.mem_writedata              (node_6_mem_writedata),                  //             .writedata
		.output_east_data           (node_6_output_east_data),               //  output_east.data
		.output_east_valid          (node_6_output_east_valid),              //             .valid
		.output_east_ready          (node_6_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_6_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_6_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_6_output_east_empty),              //             .empty
		.output_north_data          (node_6_output_north_data),              // output_north.data
		.output_north_valid         (node_6_output_north_valid),             //             .valid
		.output_north_ready         (node_6_output_north_ready),             //             .ready
		.output_north_startofpacket (node_6_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_6_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_6_output_north_empty),             //             .empty
		.output_south_data          (node_6_output_south_data),              // output_south.data
		.output_south_valid         (node_6_output_south_valid),             //             .valid
		.output_south_ready         (node_6_output_south_ready),             //             .ready
		.output_south_startofpacket (node_6_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_6_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_6_output_south_empty),             //             .empty
		.output_west_data           (node_6_output_west_data),               //  output_west.data
		.output_west_valid          (node_6_output_west_valid),              //             .valid
		.output_west_ready          (node_6_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_6_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_6_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_6_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65536 node_65536 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65537_output_west_data),            //   input_east.data
		.input_east_valid           (node_65537_output_west_valid),           //             .valid
		.input_east_ready           (node_65537_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65537_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65537_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65537_output_west_empty),           //             .empty
		.input_north_data           (node_0_output_south_data),               //  input_north.data
		.input_north_valid          (node_0_output_south_valid),              //             .valid
		.input_north_ready          (node_0_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_0_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_0_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_0_output_south_empty),              //             .empty
		.input_south_data           (node_131072_output_north_data),          //  input_south.data
		.input_south_valid          (node_131072_output_north_valid),         //             .valid
		.input_south_ready          (node_131072_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131072_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131072_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131072_output_north_empty),         //             .empty
		.input_west_data            (),                                       //   input_west.data
		.input_west_valid           (),                                       //             .valid
		.input_west_ready           (),                                       //             .ready
		.input_west_startofpacket   (),                                       //             .startofpacket
		.input_west_endofpacket     (),                                       //             .endofpacket
		.input_west_empty           (),                                       //             .empty
		.mem_address                (node_65536_mem_address),                 //          mem.address
		.mem_readdata               (node_65536_mem_readdata),                //             .readdata
		.mem_write                  (node_65536_mem_write),                   //             .write
		.mem_writedata              (node_65536_mem_writedata),               //             .writedata
		.output_east_data           (node_65536_output_east_data),            //  output_east.data
		.output_east_valid          (node_65536_output_east_valid),           //             .valid
		.output_east_ready          (node_65536_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65536_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65536_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65536_output_east_empty),           //             .empty
		.output_north_data          (node_65536_output_north_data),           // output_north.data
		.output_north_valid         (node_65536_output_north_valid),          //             .valid
		.output_north_ready         (node_65536_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65536_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65536_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65536_output_north_empty),          //             .empty
		.output_south_data          (node_65536_output_south_data),           // output_south.data
		.output_south_valid         (node_65536_output_south_valid),          //             .valid
		.output_south_ready         (node_65536_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65536_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65536_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65536_output_south_empty),          //             .empty
		.output_west_data           (node_65536_output_west_data),            //  output_west.data
		.output_west_valid          (node_65536_output_west_valid),           //             .valid
		.output_west_ready          (node_65536_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65536_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65536_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65536_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65537 node_65537 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65538_output_west_data),            //   input_east.data
		.input_east_valid           (node_65538_output_west_valid),           //             .valid
		.input_east_ready           (node_65538_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65538_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65538_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65538_output_west_empty),           //             .empty
		.input_north_data           (node_1_output_south_data),               //  input_north.data
		.input_north_valid          (node_1_output_south_valid),              //             .valid
		.input_north_ready          (node_1_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_1_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_1_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_1_output_south_empty),              //             .empty
		.input_south_data           (node_131073_output_north_data),          //  input_south.data
		.input_south_valid          (node_131073_output_north_valid),         //             .valid
		.input_south_ready          (node_131073_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131073_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131073_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131073_output_north_empty),         //             .empty
		.input_west_data            (node_65536_output_east_data),            //   input_west.data
		.input_west_valid           (node_65536_output_east_valid),           //             .valid
		.input_west_ready           (node_65536_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65536_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65536_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65536_output_east_empty),           //             .empty
		.mem_address                (node_65537_mem_address),                 //          mem.address
		.mem_readdata               (node_65537_mem_readdata),                //             .readdata
		.mem_write                  (node_65537_mem_write),                   //             .write
		.mem_writedata              (node_65537_mem_writedata),               //             .writedata
		.output_east_data           (node_65537_output_east_data),            //  output_east.data
		.output_east_valid          (node_65537_output_east_valid),           //             .valid
		.output_east_ready          (node_65537_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65537_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65537_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65537_output_east_empty),           //             .empty
		.output_north_data          (node_65537_output_north_data),           // output_north.data
		.output_north_valid         (node_65537_output_north_valid),          //             .valid
		.output_north_ready         (node_65537_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65537_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65537_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65537_output_north_empty),          //             .empty
		.output_south_data          (node_65537_output_south_data),           // output_south.data
		.output_south_valid         (node_65537_output_south_valid),          //             .valid
		.output_south_ready         (node_65537_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65537_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65537_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65537_output_south_empty),          //             .empty
		.output_west_data           (node_65537_output_west_data),            //  output_west.data
		.output_west_valid          (node_65537_output_west_valid),           //             .valid
		.output_west_ready          (node_65537_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65537_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65537_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65537_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65538 node_65538 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65539_output_west_data),            //   input_east.data
		.input_east_valid           (node_65539_output_west_valid),           //             .valid
		.input_east_ready           (node_65539_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65539_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65539_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65539_output_west_empty),           //             .empty
		.input_north_data           (node_2_output_south_data),               //  input_north.data
		.input_north_valid          (node_2_output_south_valid),              //             .valid
		.input_north_ready          (node_2_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_2_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_2_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_2_output_south_empty),              //             .empty
		.input_south_data           (node_131074_output_north_data),          //  input_south.data
		.input_south_valid          (node_131074_output_north_valid),         //             .valid
		.input_south_ready          (node_131074_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131074_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131074_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131074_output_north_empty),         //             .empty
		.input_west_data            (node_65537_output_east_data),            //   input_west.data
		.input_west_valid           (node_65537_output_east_valid),           //             .valid
		.input_west_ready           (node_65537_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65537_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65537_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65537_output_east_empty),           //             .empty
		.mem_address                (node_65538_mem_address),                 //          mem.address
		.mem_readdata               (node_65538_mem_readdata),                //             .readdata
		.mem_write                  (node_65538_mem_write),                   //             .write
		.mem_writedata              (node_65538_mem_writedata),               //             .writedata
		.output_east_data           (node_65538_output_east_data),            //  output_east.data
		.output_east_valid          (node_65538_output_east_valid),           //             .valid
		.output_east_ready          (node_65538_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65538_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65538_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65538_output_east_empty),           //             .empty
		.output_north_data          (node_65538_output_north_data),           // output_north.data
		.output_north_valid         (node_65538_output_north_valid),          //             .valid
		.output_north_ready         (node_65538_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65538_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65538_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65538_output_north_empty),          //             .empty
		.output_south_data          (node_65538_output_south_data),           // output_south.data
		.output_south_valid         (node_65538_output_south_valid),          //             .valid
		.output_south_ready         (node_65538_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65538_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65538_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65538_output_south_empty),          //             .empty
		.output_west_data           (node_65538_output_west_data),            //  output_west.data
		.output_west_valid          (node_65538_output_west_valid),           //             .valid
		.output_west_ready          (node_65538_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65538_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65538_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65538_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65539 node_65539 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65540_output_west_data),            //   input_east.data
		.input_east_valid           (node_65540_output_west_valid),           //             .valid
		.input_east_ready           (node_65540_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65540_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65540_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65540_output_west_empty),           //             .empty
		.input_north_data           (node_3_output_south_data),               //  input_north.data
		.input_north_valid          (node_3_output_south_valid),              //             .valid
		.input_north_ready          (node_3_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_3_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_3_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_3_output_south_empty),              //             .empty
		.input_south_data           (node_131075_output_north_data),          //  input_south.data
		.input_south_valid          (node_131075_output_north_valid),         //             .valid
		.input_south_ready          (node_131075_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131075_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131075_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131075_output_north_empty),         //             .empty
		.input_west_data            (node_65538_output_east_data),            //   input_west.data
		.input_west_valid           (node_65538_output_east_valid),           //             .valid
		.input_west_ready           (node_65538_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65538_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65538_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65538_output_east_empty),           //             .empty
		.mem_address                (node_65539_mem_address),                 //          mem.address
		.mem_readdata               (node_65539_mem_readdata),                //             .readdata
		.mem_write                  (node_65539_mem_write),                   //             .write
		.mem_writedata              (node_65539_mem_writedata),               //             .writedata
		.output_east_data           (node_65539_output_east_data),            //  output_east.data
		.output_east_valid          (node_65539_output_east_valid),           //             .valid
		.output_east_ready          (node_65539_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65539_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65539_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65539_output_east_empty),           //             .empty
		.output_north_data          (node_65539_output_north_data),           // output_north.data
		.output_north_valid         (node_65539_output_north_valid),          //             .valid
		.output_north_ready         (node_65539_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65539_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65539_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65539_output_north_empty),          //             .empty
		.output_south_data          (node_65539_output_south_data),           // output_south.data
		.output_south_valid         (node_65539_output_south_valid),          //             .valid
		.output_south_ready         (node_65539_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65539_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65539_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65539_output_south_empty),          //             .empty
		.output_west_data           (node_65539_output_west_data),            //  output_west.data
		.output_west_valid          (node_65539_output_west_valid),           //             .valid
		.output_west_ready          (node_65539_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65539_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65539_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65539_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65540 node_65540 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65541_output_west_data),            //   input_east.data
		.input_east_valid           (node_65541_output_west_valid),           //             .valid
		.input_east_ready           (node_65541_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65541_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65541_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65541_output_west_empty),           //             .empty
		.input_north_data           (node_4_output_south_data),               //  input_north.data
		.input_north_valid          (node_4_output_south_valid),              //             .valid
		.input_north_ready          (node_4_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_4_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_4_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_4_output_south_empty),              //             .empty
		.input_south_data           (node_131076_output_north_data),          //  input_south.data
		.input_south_valid          (node_131076_output_north_valid),         //             .valid
		.input_south_ready          (node_131076_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131076_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131076_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131076_output_north_empty),         //             .empty
		.input_west_data            (node_65539_output_east_data),            //   input_west.data
		.input_west_valid           (node_65539_output_east_valid),           //             .valid
		.input_west_ready           (node_65539_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65539_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65539_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65539_output_east_empty),           //             .empty
		.mem_address                (node_65540_mem_address),                 //          mem.address
		.mem_readdata               (node_65540_mem_readdata),                //             .readdata
		.mem_write                  (node_65540_mem_write),                   //             .write
		.mem_writedata              (node_65540_mem_writedata),               //             .writedata
		.output_east_data           (node_65540_output_east_data),            //  output_east.data
		.output_east_valid          (node_65540_output_east_valid),           //             .valid
		.output_east_ready          (node_65540_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65540_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65540_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65540_output_east_empty),           //             .empty
		.output_north_data          (node_65540_output_north_data),           // output_north.data
		.output_north_valid         (node_65540_output_north_valid),          //             .valid
		.output_north_ready         (node_65540_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65540_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65540_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65540_output_north_empty),          //             .empty
		.output_south_data          (node_65540_output_south_data),           // output_south.data
		.output_south_valid         (node_65540_output_south_valid),          //             .valid
		.output_south_ready         (node_65540_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65540_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65540_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65540_output_south_empty),          //             .empty
		.output_west_data           (node_65540_output_west_data),            //  output_west.data
		.output_west_valid          (node_65540_output_west_valid),           //             .valid
		.output_west_ready          (node_65540_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65540_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65540_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65540_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65541 node_65541 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65542_output_west_data),            //   input_east.data
		.input_east_valid           (node_65542_output_west_valid),           //             .valid
		.input_east_ready           (node_65542_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65542_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65542_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65542_output_west_empty),           //             .empty
		.input_north_data           (node_5_output_south_data),               //  input_north.data
		.input_north_valid          (node_5_output_south_valid),              //             .valid
		.input_north_ready          (node_5_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_5_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_5_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_5_output_south_empty),              //             .empty
		.input_south_data           (node_131077_output_north_data),          //  input_south.data
		.input_south_valid          (node_131077_output_north_valid),         //             .valid
		.input_south_ready          (node_131077_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131077_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131077_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131077_output_north_empty),         //             .empty
		.input_west_data            (node_65540_output_east_data),            //   input_west.data
		.input_west_valid           (node_65540_output_east_valid),           //             .valid
		.input_west_ready           (node_65540_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65540_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65540_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65540_output_east_empty),           //             .empty
		.mem_address                (node_65541_mem_address),                 //          mem.address
		.mem_readdata               (node_65541_mem_readdata),                //             .readdata
		.mem_write                  (node_65541_mem_write),                   //             .write
		.mem_writedata              (node_65541_mem_writedata),               //             .writedata
		.output_east_data           (node_65541_output_east_data),            //  output_east.data
		.output_east_valid          (node_65541_output_east_valid),           //             .valid
		.output_east_ready          (node_65541_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65541_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65541_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65541_output_east_empty),           //             .empty
		.output_north_data          (node_65541_output_north_data),           // output_north.data
		.output_north_valid         (node_65541_output_north_valid),          //             .valid
		.output_north_ready         (node_65541_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65541_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65541_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65541_output_north_empty),          //             .empty
		.output_south_data          (node_65541_output_south_data),           // output_south.data
		.output_south_valid         (node_65541_output_south_valid),          //             .valid
		.output_south_ready         (node_65541_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65541_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65541_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65541_output_south_empty),          //             .empty
		.output_west_data           (node_65541_output_west_data),            //  output_west.data
		.output_west_valid          (node_65541_output_west_valid),           //             .valid
		.output_west_ready          (node_65541_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65541_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65541_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65541_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65542 node_65542 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65543_output_west_data),            //   input_east.data
		.input_east_valid           (node_65543_output_west_valid),           //             .valid
		.input_east_ready           (node_65543_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65543_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65543_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65543_output_west_empty),           //             .empty
		.input_north_data           (node_6_output_south_data),               //  input_north.data
		.input_north_valid          (node_6_output_south_valid),              //             .valid
		.input_north_ready          (node_6_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_6_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_6_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_6_output_south_empty),              //             .empty
		.input_south_data           (node_131078_output_north_data),          //  input_south.data
		.input_south_valid          (node_131078_output_north_valid),         //             .valid
		.input_south_ready          (node_131078_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131078_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131078_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131078_output_north_empty),         //             .empty
		.input_west_data            (node_65541_output_east_data),            //   input_west.data
		.input_west_valid           (node_65541_output_east_valid),           //             .valid
		.input_west_ready           (node_65541_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65541_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65541_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65541_output_east_empty),           //             .empty
		.mem_address                (node_65542_mem_address),                 //          mem.address
		.mem_readdata               (node_65542_mem_readdata),                //             .readdata
		.mem_write                  (node_65542_mem_write),                   //             .write
		.mem_writedata              (node_65542_mem_writedata),               //             .writedata
		.output_east_data           (node_65542_output_east_data),            //  output_east.data
		.output_east_valid          (node_65542_output_east_valid),           //             .valid
		.output_east_ready          (node_65542_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65542_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65542_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65542_output_east_empty),           //             .empty
		.output_north_data          (node_65542_output_north_data),           // output_north.data
		.output_north_valid         (node_65542_output_north_valid),          //             .valid
		.output_north_ready         (node_65542_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65542_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65542_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65542_output_north_empty),          //             .empty
		.output_south_data          (node_65542_output_south_data),           // output_south.data
		.output_south_valid         (node_65542_output_south_valid),          //             .valid
		.output_south_ready         (node_65542_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65542_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65542_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65542_output_south_empty),          //             .empty
		.output_west_data           (node_65542_output_west_data),            //  output_west.data
		.output_west_valid          (node_65542_output_west_valid),           //             .valid
		.output_west_ready          (node_65542_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65542_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65542_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65542_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65543 node_65543 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (node_65544_output_west_data),            //   input_east.data
		.input_east_valid           (node_65544_output_west_valid),           //             .valid
		.input_east_ready           (node_65544_output_west_ready),           //             .ready
		.input_east_startofpacket   (node_65544_output_west_startofpacket),   //             .startofpacket
		.input_east_endofpacket     (node_65544_output_west_endofpacket),     //             .endofpacket
		.input_east_empty           (node_65544_output_west_empty),           //             .empty
		.input_north_data           (node_7_output_south_data),               //  input_north.data
		.input_north_valid          (node_7_output_south_valid),              //             .valid
		.input_north_ready          (node_7_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_7_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_7_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_7_output_south_empty),              //             .empty
		.input_south_data           (node_131079_output_north_data),          //  input_south.data
		.input_south_valid          (node_131079_output_north_valid),         //             .valid
		.input_south_ready          (node_131079_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131079_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131079_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131079_output_north_empty),         //             .empty
		.input_west_data            (node_65542_output_east_data),            //   input_west.data
		.input_west_valid           (node_65542_output_east_valid),           //             .valid
		.input_west_ready           (node_65542_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65542_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65542_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65542_output_east_empty),           //             .empty
		.mem_address                (node_65543_mem_address),                 //          mem.address
		.mem_readdata               (node_65543_mem_readdata),                //             .readdata
		.mem_write                  (node_65543_mem_write),                   //             .write
		.mem_writedata              (node_65543_mem_writedata),               //             .writedata
		.output_east_data           (node_65543_output_east_data),            //  output_east.data
		.output_east_valid          (node_65543_output_east_valid),           //             .valid
		.output_east_ready          (node_65543_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65543_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65543_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65543_output_east_empty),           //             .empty
		.output_north_data          (node_65543_output_north_data),           // output_north.data
		.output_north_valid         (node_65543_output_north_valid),          //             .valid
		.output_north_ready         (node_65543_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65543_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65543_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65543_output_north_empty),          //             .empty
		.output_south_data          (node_65543_output_south_data),           // output_south.data
		.output_south_valid         (node_65543_output_south_valid),          //             .valid
		.output_south_ready         (node_65543_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65543_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65543_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65543_output_south_empty),          //             .empty
		.output_west_data           (node_65543_output_west_data),            //  output_west.data
		.output_west_valid          (node_65543_output_west_valid),           //             .valid
		.output_west_ready          (node_65543_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65543_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65543_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65543_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_65544 node_65544 (
		.clk_clk                    (clk_clk),                                //          clk.clk
		.input_east_data            (),                                       //   input_east.data
		.input_east_valid           (),                                       //             .valid
		.input_east_ready           (),                                       //             .ready
		.input_east_startofpacket   (),                                       //             .startofpacket
		.input_east_endofpacket     (),                                       //             .endofpacket
		.input_east_empty           (),                                       //             .empty
		.input_north_data           (node_8_output_south_data),               //  input_north.data
		.input_north_valid          (node_8_output_south_valid),              //             .valid
		.input_north_ready          (node_8_output_south_ready),              //             .ready
		.input_north_startofpacket  (node_8_output_south_startofpacket),      //             .startofpacket
		.input_north_endofpacket    (node_8_output_south_endofpacket),        //             .endofpacket
		.input_north_empty          (node_8_output_south_empty),              //             .empty
		.input_south_data           (node_131080_output_north_data),          //  input_south.data
		.input_south_valid          (node_131080_output_north_valid),         //             .valid
		.input_south_ready          (node_131080_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_131080_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_131080_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_131080_output_north_empty),         //             .empty
		.input_west_data            (node_65543_output_east_data),            //   input_west.data
		.input_west_valid           (node_65543_output_east_valid),           //             .valid
		.input_west_ready           (node_65543_output_east_ready),           //             .ready
		.input_west_startofpacket   (node_65543_output_east_startofpacket),   //             .startofpacket
		.input_west_endofpacket     (node_65543_output_east_endofpacket),     //             .endofpacket
		.input_west_empty           (node_65543_output_east_empty),           //             .empty
		.mem_address                (node_65544_mem_address),                 //          mem.address
		.mem_readdata               (node_65544_mem_readdata),                //             .readdata
		.mem_write                  (node_65544_mem_write),                   //             .write
		.mem_writedata              (node_65544_mem_writedata),               //             .writedata
		.output_east_data           (node_65544_output_east_data),            //  output_east.data
		.output_east_valid          (node_65544_output_east_valid),           //             .valid
		.output_east_ready          (node_65544_output_east_ready),           //             .ready
		.output_east_startofpacket  (node_65544_output_east_startofpacket),   //             .startofpacket
		.output_east_endofpacket    (node_65544_output_east_endofpacket),     //             .endofpacket
		.output_east_empty          (node_65544_output_east_empty),           //             .empty
		.output_north_data          (node_65544_output_north_data),           // output_north.data
		.output_north_valid         (node_65544_output_north_valid),          //             .valid
		.output_north_ready         (node_65544_output_north_ready),          //             .ready
		.output_north_startofpacket (node_65544_output_north_startofpacket),  //             .startofpacket
		.output_north_endofpacket   (node_65544_output_north_endofpacket),    //             .endofpacket
		.output_north_empty         (node_65544_output_north_empty),          //             .empty
		.output_south_data          (node_65544_output_south_data),           // output_south.data
		.output_south_valid         (node_65544_output_south_valid),          //             .valid
		.output_south_ready         (node_65544_output_south_ready),          //             .ready
		.output_south_startofpacket (node_65544_output_south_startofpacket),  //             .startofpacket
		.output_south_endofpacket   (node_65544_output_south_endofpacket),    //             .endofpacket
		.output_south_empty         (node_65544_output_south_empty),          //             .empty
		.output_west_data           (node_65544_output_west_data),            //  output_west.data
		.output_west_valid          (node_65544_output_west_valid),           //             .valid
		.output_west_ready          (node_65544_output_west_ready),           //             .ready
		.output_west_startofpacket  (node_65544_output_west_startofpacket),   //             .startofpacket
		.output_west_endofpacket    (node_65544_output_west_endofpacket),     //             .endofpacket
		.output_west_empty          (node_65544_output_west_empty),           //             .empty
		.reset_reset_n              (reset_reset_n)                           //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_7 node_7 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (node_8_output_west_data),               //   input_east.data
		.input_east_valid           (node_8_output_west_valid),              //             .valid
		.input_east_ready           (node_8_output_west_ready),              //             .ready
		.input_east_startofpacket   (node_8_output_west_startofpacket),      //             .startofpacket
		.input_east_endofpacket     (node_8_output_west_endofpacket),        //             .endofpacket
		.input_east_empty           (node_8_output_west_empty),              //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65543_output_north_data),          //  input_south.data
		.input_south_valid          (node_65543_output_north_valid),         //             .valid
		.input_south_ready          (node_65543_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65543_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65543_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65543_output_north_empty),         //             .empty
		.input_west_data            (node_6_output_east_data),               //   input_west.data
		.input_west_valid           (node_6_output_east_valid),              //             .valid
		.input_west_ready           (node_6_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_6_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_6_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_6_output_east_empty),              //             .empty
		.mem_address                (node_7_mem_address),                    //          mem.address
		.mem_readdata               (node_7_mem_readdata),                   //             .readdata
		.mem_write                  (node_7_mem_write),                      //             .write
		.mem_writedata              (node_7_mem_writedata),                  //             .writedata
		.output_east_data           (node_7_output_east_data),               //  output_east.data
		.output_east_valid          (node_7_output_east_valid),              //             .valid
		.output_east_ready          (node_7_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_7_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_7_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_7_output_east_empty),              //             .empty
		.output_north_data          (node_7_output_north_data),              // output_north.data
		.output_north_valid         (node_7_output_north_valid),             //             .valid
		.output_north_ready         (node_7_output_north_ready),             //             .ready
		.output_north_startofpacket (node_7_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_7_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_7_output_north_empty),             //             .empty
		.output_south_data          (node_7_output_south_data),              // output_south.data
		.output_south_valid         (node_7_output_south_valid),             //             .valid
		.output_south_ready         (node_7_output_south_ready),             //             .ready
		.output_south_startofpacket (node_7_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_7_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_7_output_south_empty),             //             .empty
		.output_west_data           (node_7_output_west_data),               //  output_west.data
		.output_west_valid          (node_7_output_west_valid),              //             .valid
		.output_west_ready          (node_7_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_7_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_7_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_7_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_system_rtl_gals_test_version_node_8 node_8 (
		.clk_clk                    (clk_clk),                               //          clk.clk
		.input_east_data            (),                                      //   input_east.data
		.input_east_valid           (),                                      //             .valid
		.input_east_ready           (),                                      //             .ready
		.input_east_startofpacket   (),                                      //             .startofpacket
		.input_east_endofpacket     (),                                      //             .endofpacket
		.input_east_empty           (),                                      //             .empty
		.input_north_data           (),                                      //  input_north.data
		.input_north_valid          (),                                      //             .valid
		.input_north_ready          (),                                      //             .ready
		.input_north_startofpacket  (),                                      //             .startofpacket
		.input_north_endofpacket    (),                                      //             .endofpacket
		.input_north_empty          (),                                      //             .empty
		.input_south_data           (node_65544_output_north_data),          //  input_south.data
		.input_south_valid          (node_65544_output_north_valid),         //             .valid
		.input_south_ready          (node_65544_output_north_ready),         //             .ready
		.input_south_startofpacket  (node_65544_output_north_startofpacket), //             .startofpacket
		.input_south_endofpacket    (node_65544_output_north_endofpacket),   //             .endofpacket
		.input_south_empty          (node_65544_output_north_empty),         //             .empty
		.input_west_data            (node_7_output_east_data),               //   input_west.data
		.input_west_valid           (node_7_output_east_valid),              //             .valid
		.input_west_ready           (node_7_output_east_ready),              //             .ready
		.input_west_startofpacket   (node_7_output_east_startofpacket),      //             .startofpacket
		.input_west_endofpacket     (node_7_output_east_endofpacket),        //             .endofpacket
		.input_west_empty           (node_7_output_east_empty),              //             .empty
		.mem_address                (node_8_mem_address),                    //          mem.address
		.mem_readdata               (node_8_mem_readdata),                   //             .readdata
		.mem_write                  (node_8_mem_write),                      //             .write
		.mem_writedata              (node_8_mem_writedata),                  //             .writedata
		.output_east_data           (node_8_output_east_data),               //  output_east.data
		.output_east_valid          (node_8_output_east_valid),              //             .valid
		.output_east_ready          (node_8_output_east_ready),              //             .ready
		.output_east_startofpacket  (node_8_output_east_startofpacket),      //             .startofpacket
		.output_east_endofpacket    (node_8_output_east_endofpacket),        //             .endofpacket
		.output_east_empty          (node_8_output_east_empty),              //             .empty
		.output_north_data          (node_8_output_north_data),              // output_north.data
		.output_north_valid         (node_8_output_north_valid),             //             .valid
		.output_north_ready         (node_8_output_north_ready),             //             .ready
		.output_north_startofpacket (node_8_output_north_startofpacket),     //             .startofpacket
		.output_north_endofpacket   (node_8_output_north_endofpacket),       //             .endofpacket
		.output_north_empty         (node_8_output_north_empty),             //             .empty
		.output_south_data          (node_8_output_south_data),              // output_south.data
		.output_south_valid         (node_8_output_south_valid),             //             .valid
		.output_south_ready         (node_8_output_south_ready),             //             .ready
		.output_south_startofpacket (node_8_output_south_startofpacket),     //             .startofpacket
		.output_south_endofpacket   (node_8_output_south_endofpacket),       //             .endofpacket
		.output_south_empty         (node_8_output_south_empty),             //             .empty
		.output_west_data           (node_8_output_west_data),               //  output_west.data
		.output_west_valid          (node_8_output_west_valid),              //             .valid
		.output_west_ready          (node_8_output_west_ready),              //             .ready
		.output_west_startofpacket  (node_8_output_west_startofpacket),      //             .startofpacket
		.output_west_endofpacket    (node_8_output_west_endofpacket),        //             .endofpacket
		.output_west_empty          (node_8_output_west_empty),              //             .empty
		.reset_reset_n              (reset_reset_n)                          //        reset.reset_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_east_0 (
		.reset_n       (~rst_controller_reset_out_reset),  //  reset.reset_n
		.clk           (clk_clk),                          //  clock.clk
		.data          (node_8_output_east_data),          //     s1.data
		.empty         (node_8_output_east_empty),         //       .empty
		.endofpacket   (node_8_output_east_endofpacket),   //       .endofpacket
		.ready         (node_8_output_east_ready),         //       .ready
		.startofpacket (node_8_output_east_startofpacket), //       .startofpacket
		.valid         (node_8_output_east_valid),         //       .valid
		.readdata      (),                                 // status.readdata
		.address       (),                                 //       .address
		.read_n        ()                                  //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_east_1 (
		.reset_n       (~rst_controller_reset_out_reset),      //  reset.reset_n
		.clk           (clk_clk),                              //  clock.clk
		.data          (node_65544_output_east_data),          //     s1.data
		.empty         (node_65544_output_east_empty),         //       .empty
		.endofpacket   (node_65544_output_east_endofpacket),   //       .endofpacket
		.ready         (node_65544_output_east_ready),         //       .ready
		.startofpacket (node_65544_output_east_startofpacket), //       .startofpacket
		.valid         (node_65544_output_east_valid),         //       .valid
		.readdata      (),                                     // status.readdata
		.address       (),                                     //       .address
		.read_n        ()                                      //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_east_2 (
		.reset_n       (~rst_controller_reset_out_reset),       //  reset.reset_n
		.clk           (clk_clk),                               //  clock.clk
		.data          (node_131080_output_east_data),          //     s1.data
		.empty         (node_131080_output_east_empty),         //       .empty
		.endofpacket   (node_131080_output_east_endofpacket),   //       .endofpacket
		.ready         (node_131080_output_east_ready),         //       .ready
		.startofpacket (node_131080_output_east_startofpacket), //       .startofpacket
		.valid         (node_131080_output_east_valid),         //       .valid
		.readdata      (),                                      // status.readdata
		.address       (),                                      //       .address
		.read_n        ()                                       //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_0 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_0_output_north_data),          //     s1.data
		.empty         (node_0_output_north_empty),         //       .empty
		.endofpacket   (node_0_output_north_endofpacket),   //       .endofpacket
		.ready         (node_0_output_north_ready),         //       .ready
		.startofpacket (node_0_output_north_startofpacket), //       .startofpacket
		.valid         (node_0_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_1 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_1_output_north_data),          //     s1.data
		.empty         (node_1_output_north_empty),         //       .empty
		.endofpacket   (node_1_output_north_endofpacket),   //       .endofpacket
		.ready         (node_1_output_north_ready),         //       .ready
		.startofpacket (node_1_output_north_startofpacket), //       .startofpacket
		.valid         (node_1_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_2 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_2_output_north_data),          //     s1.data
		.empty         (node_2_output_north_empty),         //       .empty
		.endofpacket   (node_2_output_north_endofpacket),   //       .endofpacket
		.ready         (node_2_output_north_ready),         //       .ready
		.startofpacket (node_2_output_north_startofpacket), //       .startofpacket
		.valid         (node_2_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_3 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_3_output_north_data),          //     s1.data
		.empty         (node_3_output_north_empty),         //       .empty
		.endofpacket   (node_3_output_north_endofpacket),   //       .endofpacket
		.ready         (node_3_output_north_ready),         //       .ready
		.startofpacket (node_3_output_north_startofpacket), //       .startofpacket
		.valid         (node_3_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_4 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_4_output_north_data),          //     s1.data
		.empty         (node_4_output_north_empty),         //       .empty
		.endofpacket   (node_4_output_north_endofpacket),   //       .endofpacket
		.ready         (node_4_output_north_ready),         //       .ready
		.startofpacket (node_4_output_north_startofpacket), //       .startofpacket
		.valid         (node_4_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_5 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_5_output_north_data),          //     s1.data
		.empty         (node_5_output_north_empty),         //       .empty
		.endofpacket   (node_5_output_north_endofpacket),   //       .endofpacket
		.ready         (node_5_output_north_ready),         //       .ready
		.startofpacket (node_5_output_north_startofpacket), //       .startofpacket
		.valid         (node_5_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_6 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_6_output_north_data),          //     s1.data
		.empty         (node_6_output_north_empty),         //       .empty
		.endofpacket   (node_6_output_north_endofpacket),   //       .endofpacket
		.ready         (node_6_output_north_ready),         //       .ready
		.startofpacket (node_6_output_north_startofpacket), //       .startofpacket
		.valid         (node_6_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_7 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_7_output_north_data),          //     s1.data
		.empty         (node_7_output_north_empty),         //       .empty
		.endofpacket   (node_7_output_north_endofpacket),   //       .endofpacket
		.ready         (node_7_output_north_ready),         //       .ready
		.startofpacket (node_7_output_north_startofpacket), //       .startofpacket
		.valid         (node_7_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_north_8 (
		.reset_n       (~rst_controller_reset_out_reset),   //  reset.reset_n
		.clk           (clk_clk),                           //  clock.clk
		.data          (node_8_output_north_data),          //     s1.data
		.empty         (node_8_output_north_empty),         //       .empty
		.endofpacket   (node_8_output_north_endofpacket),   //       .endofpacket
		.ready         (node_8_output_north_ready),         //       .ready
		.startofpacket (node_8_output_north_startofpacket), //       .startofpacket
		.valid         (node_8_output_north_valid),         //       .valid
		.readdata      (),                                  // status.readdata
		.address       (),                                  //       .address
		.read_n        ()                                   //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_0 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131072_output_south_data),          //     s1.data
		.empty         (node_131072_output_south_empty),         //       .empty
		.endofpacket   (node_131072_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131072_output_south_ready),         //       .ready
		.startofpacket (node_131072_output_south_startofpacket), //       .startofpacket
		.valid         (node_131072_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_1 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131073_output_south_data),          //     s1.data
		.empty         (node_131073_output_south_empty),         //       .empty
		.endofpacket   (node_131073_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131073_output_south_ready),         //       .ready
		.startofpacket (node_131073_output_south_startofpacket), //       .startofpacket
		.valid         (node_131073_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_2 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131074_output_south_data),          //     s1.data
		.empty         (node_131074_output_south_empty),         //       .empty
		.endofpacket   (node_131074_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131074_output_south_ready),         //       .ready
		.startofpacket (node_131074_output_south_startofpacket), //       .startofpacket
		.valid         (node_131074_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_3 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131075_output_south_data),          //     s1.data
		.empty         (node_131075_output_south_empty),         //       .empty
		.endofpacket   (node_131075_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131075_output_south_ready),         //       .ready
		.startofpacket (node_131075_output_south_startofpacket), //       .startofpacket
		.valid         (node_131075_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_4 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131076_output_south_data),          //     s1.data
		.empty         (node_131076_output_south_empty),         //       .empty
		.endofpacket   (node_131076_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131076_output_south_ready),         //       .ready
		.startofpacket (node_131076_output_south_startofpacket), //       .startofpacket
		.valid         (node_131076_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_5 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131077_output_south_data),          //     s1.data
		.empty         (node_131077_output_south_empty),         //       .empty
		.endofpacket   (node_131077_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131077_output_south_ready),         //       .ready
		.startofpacket (node_131077_output_south_startofpacket), //       .startofpacket
		.valid         (node_131077_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_6 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131078_output_south_data),          //     s1.data
		.empty         (node_131078_output_south_empty),         //       .empty
		.endofpacket   (node_131078_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131078_output_south_ready),         //       .ready
		.startofpacket (node_131078_output_south_startofpacket), //       .startofpacket
		.valid         (node_131078_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_7 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131079_output_south_data),          //     s1.data
		.empty         (node_131079_output_south_empty),         //       .empty
		.endofpacket   (node_131079_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131079_output_south_ready),         //       .ready
		.startofpacket (node_131079_output_south_startofpacket), //       .startofpacket
		.valid         (node_131079_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_south_8 (
		.reset_n       (~rst_controller_reset_out_reset),        //  reset.reset_n
		.clk           (clk_clk),                                //  clock.clk
		.data          (node_131080_output_south_data),          //     s1.data
		.empty         (node_131080_output_south_empty),         //       .empty
		.endofpacket   (node_131080_output_south_endofpacket),   //       .endofpacket
		.ready         (node_131080_output_south_ready),         //       .ready
		.startofpacket (node_131080_output_south_startofpacket), //       .startofpacket
		.valid         (node_131080_output_south_valid),         //       .valid
		.readdata      (),                                       // status.readdata
		.address       (),                                       //       .address
		.read_n        ()                                        //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_west_0 (
		.reset_n       (~rst_controller_reset_out_reset),  //  reset.reset_n
		.clk           (clk_clk),                          //  clock.clk
		.data          (node_0_output_west_data),          //     s1.data
		.empty         (node_0_output_west_empty),         //       .empty
		.endofpacket   (node_0_output_west_endofpacket),   //       .endofpacket
		.ready         (node_0_output_west_ready),         //       .ready
		.startofpacket (node_0_output_west_startofpacket), //       .startofpacket
		.valid         (node_0_output_west_valid),         //       .valid
		.readdata      (),                                 // status.readdata
		.address       (),                                 //       .address
		.read_n        ()                                  //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_west_1 (
		.reset_n       (~rst_controller_reset_out_reset),      //  reset.reset_n
		.clk           (clk_clk),                              //  clock.clk
		.data          (node_65536_output_west_data),          //     s1.data
		.empty         (node_65536_output_west_empty),         //       .empty
		.endofpacket   (node_65536_output_west_endofpacket),   //       .endofpacket
		.ready         (node_65536_output_west_ready),         //       .ready
		.startofpacket (node_65536_output_west_startofpacket), //       .startofpacket
		.valid         (node_65536_output_west_valid),         //       .valid
		.readdata      (),                                     // status.readdata
		.address       (),                                     //       .address
		.read_n        ()                                      //       .read_n
	);

	dircc_avalon_st_terminal_inst #(
		.DATA_WIDTH (32)
	) terminal_west_2 (
		.reset_n       (~rst_controller_reset_out_reset),       //  reset.reset_n
		.clk           (clk_clk),                               //  clock.clk
		.data          (node_131072_output_west_data),          //     s1.data
		.empty         (node_131072_output_west_empty),         //       .empty
		.endofpacket   (node_131072_output_west_endofpacket),   //       .endofpacket
		.ready         (node_131072_output_west_ready),         //       .ready
		.startofpacket (node_131072_output_west_startofpacket), //       .startofpacket
		.valid         (node_131072_output_west_valid),         //       .valid
		.readdata      (),                                      // status.readdata
		.address       (),                                      //       .address
		.read_n        ()                                       //       .read_n
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
