// poets_routing.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module poets_routing (
		input  wire        clk_clk,                    //          clk.clk
		input  wire [31:0] input_east_data,            //   input_east.data
		input  wire        input_east_valid,           //             .valid
		output wire        input_east_ready,           //             .ready
		input  wire        input_east_startofpacket,   //             .startofpacket
		input  wire        input_east_endofpacket,     //             .endofpacket
		input  wire [1:0]  input_east_empty,           //             .empty
		input  wire [31:0] input_north_data,           //  input_north.data
		input  wire        input_north_valid,          //             .valid
		output wire        input_north_ready,          //             .ready
		input  wire        input_north_startofpacket,  //             .startofpacket
		input  wire        input_north_endofpacket,    //             .endofpacket
		input  wire [1:0]  input_north_empty,          //             .empty
		input  wire [31:0] input_poets_data,           //  input_poets.data
		input  wire        input_poets_valid,          //             .valid
		output wire        input_poets_ready,          //             .ready
		input  wire        input_poets_startofpacket,  //             .startofpacket
		input  wire        input_poets_endofpacket,    //             .endofpacket
		input  wire [1:0]  input_poets_empty,          //             .empty
		input  wire [31:0] input_south_data,           //  input_south.data
		input  wire        input_south_valid,          //             .valid
		output wire        input_south_ready,          //             .ready
		input  wire        input_south_startofpacket,  //             .startofpacket
		input  wire        input_south_endofpacket,    //             .endofpacket
		input  wire [1:0]  input_south_empty,          //             .empty
		input  wire [31:0] input_west_data,            //   input_west.data
		input  wire        input_west_valid,           //             .valid
		output wire        input_west_ready,           //             .ready
		input  wire        input_west_startofpacket,   //             .startofpacket
		input  wire        input_west_endofpacket,     //             .endofpacket
		input  wire [1:0]  input_west_empty,           //             .empty
		output wire [31:0] output_east_data,           //  output_east.data
		output wire        output_east_valid,          //             .valid
		input  wire        output_east_ready,          //             .ready
		output wire        output_east_startofpacket,  //             .startofpacket
		output wire        output_east_endofpacket,    //             .endofpacket
		output wire [1:0]  output_east_empty,          //             .empty
		output wire [31:0] output_north_data,          // output_north.data
		output wire        output_north_valid,         //             .valid
		input  wire        output_north_ready,         //             .ready
		output wire        output_north_startofpacket, //             .startofpacket
		output wire        output_north_endofpacket,   //             .endofpacket
		output wire [1:0]  output_north_empty,         //             .empty
		output wire [31:0] output_poets_data,          // output_poets.data
		output wire        output_poets_valid,         //             .valid
		input  wire        output_poets_ready,         //             .ready
		output wire        output_poets_startofpacket, //             .startofpacket
		output wire        output_poets_endofpacket,   //             .endofpacket
		output wire [1:0]  output_poets_empty,         //             .empty
		output wire [31:0] output_south_data,          // output_south.data
		output wire        output_south_valid,         //             .valid
		input  wire        output_south_ready,         //             .ready
		output wire        output_south_startofpacket, //             .startofpacket
		output wire        output_south_endofpacket,   //             .endofpacket
		output wire [1:0]  output_south_empty,         //             .empty
		output wire [31:0] output_west_data,           //  output_west.data
		output wire        output_west_valid,          //             .valid
		input  wire        output_west_ready,          //             .ready
		output wire        output_west_startofpacket,  //             .startofpacket
		output wire        output_west_endofpacket,    //             .endofpacket
		output wire [1:0]  output_west_empty,          //             .empty
		input  wire        reset_reset_n               //        reset.reset_n
	);

	wire         input_mux_out_valid;            // input_mux:out_valid -> output_demux:in_valid
	wire  [31:0] input_mux_out_data;             // input_mux:out_data -> output_demux:in_data
	wire         input_mux_out_ready;            // output_demux:in_ready -> input_mux:out_ready
	wire   [2:0] input_mux_out_channel;          // input_mux:out_channel -> output_demux:in_channel
	wire         input_mux_out_startofpacket;    // input_mux:out_startofpacket -> output_demux:in_startofpacket
	wire         input_mux_out_endofpacket;      // input_mux:out_endofpacket -> output_demux:in_endofpacket
	wire   [1:0] input_mux_out_empty;            // input_mux:out_empty -> output_demux:in_empty
	wire         input_fifo_4_out_valid;         // input_fifo_4:out_valid -> input_mux:in1_valid
	wire  [31:0] input_fifo_4_out_data;          // input_fifo_4:out_data -> input_mux:in1_data
	wire         input_fifo_4_out_ready;         // input_mux:in1_ready -> input_fifo_4:out_ready
	wire         input_fifo_4_out_startofpacket; // input_fifo_4:out_startofpacket -> input_mux:in1_startofpacket
	wire         input_fifo_4_out_endofpacket;   // input_fifo_4:out_endofpacket -> input_mux:in1_endofpacket
	wire   [1:0] input_fifo_4_out_empty;         // input_fifo_4:out_empty -> input_mux:in1_empty
	wire         input_fifo_2_out_valid;         // input_fifo_2:out_valid -> input_mux:in2_valid
	wire  [31:0] input_fifo_2_out_data;          // input_fifo_2:out_data -> input_mux:in2_data
	wire         input_fifo_2_out_ready;         // input_mux:in2_ready -> input_fifo_2:out_ready
	wire         input_fifo_2_out_startofpacket; // input_fifo_2:out_startofpacket -> input_mux:in2_startofpacket
	wire         input_fifo_2_out_endofpacket;   // input_fifo_2:out_endofpacket -> input_mux:in2_endofpacket
	wire   [1:0] input_fifo_2_out_empty;         // input_fifo_2:out_empty -> input_mux:in2_empty
	wire         input_fifo_1_out_valid;         // input_fifo_1:out_valid -> input_mux:in3_valid
	wire  [31:0] input_fifo_1_out_data;          // input_fifo_1:out_data -> input_mux:in3_data
	wire         input_fifo_1_out_ready;         // input_mux:in3_ready -> input_fifo_1:out_ready
	wire         input_fifo_1_out_startofpacket; // input_fifo_1:out_startofpacket -> input_mux:in3_startofpacket
	wire         input_fifo_1_out_endofpacket;   // input_fifo_1:out_endofpacket -> input_mux:in3_endofpacket
	wire   [1:0] input_fifo_1_out_empty;         // input_fifo_1:out_empty -> input_mux:in3_empty
	wire         input_fifo_0_out_valid;         // input_fifo_0:out_valid -> input_mux:in4_valid
	wire  [31:0] input_fifo_0_out_data;          // input_fifo_0:out_data -> input_mux:in4_data
	wire         input_fifo_0_out_ready;         // input_mux:in4_ready -> input_fifo_0:out_ready
	wire         input_fifo_0_out_startofpacket; // input_fifo_0:out_startofpacket -> input_mux:in4_startofpacket
	wire         input_fifo_0_out_endofpacket;   // input_fifo_0:out_endofpacket -> input_mux:in4_endofpacket
	wire   [1:0] input_fifo_0_out_empty;         // input_fifo_0:out_empty -> input_mux:in4_empty
	wire         rst_controller_reset_out_reset; // rst_controller:reset_out -> [input_fifo_0:reset, input_fifo_1:reset, input_fifo_2:reset, input_fifo_4:reset, input_mux:reset_n, output_demux:reset_n]

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (4),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_fifo_0 (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (input_north_data),                     //        in.data
		.in_valid          (input_north_valid),                    //          .valid
		.in_ready          (input_north_ready),                    //          .ready
		.in_startofpacket  (input_north_startofpacket),            //          .startofpacket
		.in_endofpacket    (input_north_endofpacket),              //          .endofpacket
		.in_empty          (input_north_empty),                    //          .empty
		.out_data          (input_fifo_0_out_data),                //       out.data
		.out_valid         (input_fifo_0_out_valid),               //          .valid
		.out_ready         (input_fifo_0_out_ready),               //          .ready
		.out_startofpacket (input_fifo_0_out_startofpacket),       //          .startofpacket
		.out_endofpacket   (input_fifo_0_out_endofpacket),         //          .endofpacket
		.out_empty         (input_fifo_0_out_empty),               //          .empty
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (4),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_fifo_1 (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (input_west_data),                      //        in.data
		.in_valid          (input_west_valid),                     //          .valid
		.in_ready          (input_west_ready),                     //          .ready
		.in_startofpacket  (input_west_startofpacket),             //          .startofpacket
		.in_endofpacket    (input_west_endofpacket),               //          .endofpacket
		.in_empty          (input_west_empty),                     //          .empty
		.out_data          (input_fifo_1_out_data),                //       out.data
		.out_valid         (input_fifo_1_out_valid),               //          .valid
		.out_ready         (input_fifo_1_out_ready),               //          .ready
		.out_startofpacket (input_fifo_1_out_startofpacket),       //          .startofpacket
		.out_endofpacket   (input_fifo_1_out_endofpacket),         //          .endofpacket
		.out_empty         (input_fifo_1_out_empty),               //          .empty
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (4),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_fifo_2 (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (input_east_data),                      //        in.data
		.in_valid          (input_east_valid),                     //          .valid
		.in_ready          (input_east_ready),                     //          .ready
		.in_startofpacket  (input_east_startofpacket),             //          .startofpacket
		.in_endofpacket    (input_east_endofpacket),               //          .endofpacket
		.in_empty          (input_east_empty),                     //          .empty
		.out_data          (input_fifo_2_out_data),                //       out.data
		.out_valid         (input_fifo_2_out_valid),               //          .valid
		.out_ready         (input_fifo_2_out_ready),               //          .ready
		.out_startofpacket (input_fifo_2_out_startofpacket),       //          .startofpacket
		.out_endofpacket   (input_fifo_2_out_endofpacket),         //          .endofpacket
		.out_empty         (input_fifo_2_out_empty),               //          .empty
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (4),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (16),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_fifo_4 (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (input_south_data),                     //        in.data
		.in_valid          (input_south_valid),                    //          .valid
		.in_ready          (input_south_ready),                    //          .ready
		.in_startofpacket  (input_south_startofpacket),            //          .startofpacket
		.in_endofpacket    (input_south_endofpacket),              //          .endofpacket
		.in_empty          (input_south_empty),                    //          .empty
		.out_data          (input_fifo_4_out_data),                //       out.data
		.out_valid         (input_fifo_4_out_valid),               //          .valid
		.out_ready         (input_fifo_4_out_ready),               //          .ready
		.out_startofpacket (input_fifo_4_out_startofpacket),       //          .startofpacket
		.out_endofpacket   (input_fifo_4_out_endofpacket),         //          .endofpacket
		.out_empty         (input_fifo_4_out_empty),               //          .empty
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	poets_routing_input_mux input_mux (
		.clk               (clk_clk),                         //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset), // reset.reset_n
		.out_data          (input_mux_out_data),              //   out.data
		.out_valid         (input_mux_out_valid),             //      .valid
		.out_ready         (input_mux_out_ready),             //      .ready
		.out_startofpacket (input_mux_out_startofpacket),     //      .startofpacket
		.out_endofpacket   (input_mux_out_endofpacket),       //      .endofpacket
		.out_empty         (input_mux_out_empty),             //      .empty
		.out_channel       (input_mux_out_channel),           //      .channel
		.in0_data          (input_poets_data),                //   in0.data
		.in0_valid         (input_poets_valid),               //      .valid
		.in0_ready         (input_poets_ready),               //      .ready
		.in0_startofpacket (input_poets_startofpacket),       //      .startofpacket
		.in0_endofpacket   (input_poets_endofpacket),         //      .endofpacket
		.in0_empty         (input_poets_empty),               //      .empty
		.in1_data          (input_fifo_4_out_data),           //   in1.data
		.in1_valid         (input_fifo_4_out_valid),          //      .valid
		.in1_ready         (input_fifo_4_out_ready),          //      .ready
		.in1_startofpacket (input_fifo_4_out_startofpacket),  //      .startofpacket
		.in1_endofpacket   (input_fifo_4_out_endofpacket),    //      .endofpacket
		.in1_empty         (input_fifo_4_out_empty),          //      .empty
		.in2_data          (input_fifo_2_out_data),           //   in2.data
		.in2_valid         (input_fifo_2_out_valid),          //      .valid
		.in2_ready         (input_fifo_2_out_ready),          //      .ready
		.in2_startofpacket (input_fifo_2_out_startofpacket),  //      .startofpacket
		.in2_endofpacket   (input_fifo_2_out_endofpacket),    //      .endofpacket
		.in2_empty         (input_fifo_2_out_empty),          //      .empty
		.in3_data          (input_fifo_1_out_data),           //   in3.data
		.in3_valid         (input_fifo_1_out_valid),          //      .valid
		.in3_ready         (input_fifo_1_out_ready),          //      .ready
		.in3_startofpacket (input_fifo_1_out_startofpacket),  //      .startofpacket
		.in3_endofpacket   (input_fifo_1_out_endofpacket),    //      .endofpacket
		.in3_empty         (input_fifo_1_out_empty),          //      .empty
		.in4_data          (input_fifo_0_out_data),           //   in4.data
		.in4_valid         (input_fifo_0_out_valid),          //      .valid
		.in4_ready         (input_fifo_0_out_ready),          //      .ready
		.in4_startofpacket (input_fifo_0_out_startofpacket),  //      .startofpacket
		.in4_endofpacket   (input_fifo_0_out_endofpacket),    //      .endofpacket
		.in4_empty         (input_fifo_0_out_empty)           //      .empty
	);

	poets_routing_output_demux output_demux (
		.clk                (clk_clk),                         //   clk.clk
		.reset_n            (~rst_controller_reset_out_reset), // reset.reset_n
		.in_data            (input_mux_out_data),              //    in.data
		.in_valid           (input_mux_out_valid),             //      .valid
		.in_ready           (input_mux_out_ready),             //      .ready
		.in_startofpacket   (input_mux_out_startofpacket),     //      .startofpacket
		.in_endofpacket     (input_mux_out_endofpacket),       //      .endofpacket
		.in_empty           (input_mux_out_empty),             //      .empty
		.in_channel         (input_mux_out_channel),           //      .channel
		.out0_data          (output_poets_data),               //  out0.data
		.out0_valid         (output_poets_valid),              //      .valid
		.out0_ready         (output_poets_ready),              //      .ready
		.out0_startofpacket (output_poets_startofpacket),      //      .startofpacket
		.out0_endofpacket   (output_poets_endofpacket),        //      .endofpacket
		.out0_empty         (output_poets_empty),              //      .empty
		.out1_data          (output_north_data),               //  out1.data
		.out1_valid         (output_north_valid),              //      .valid
		.out1_ready         (output_north_ready),              //      .ready
		.out1_startofpacket (output_north_startofpacket),      //      .startofpacket
		.out1_endofpacket   (output_north_endofpacket),        //      .endofpacket
		.out1_empty         (output_north_empty),              //      .empty
		.out2_data          (output_west_data),                //  out2.data
		.out2_valid         (output_west_valid),               //      .valid
		.out2_ready         (output_west_ready),               //      .ready
		.out2_startofpacket (output_west_startofpacket),       //      .startofpacket
		.out2_endofpacket   (output_west_endofpacket),         //      .endofpacket
		.out2_empty         (output_west_empty),               //      .empty
		.out3_data          (output_south_data),               //  out3.data
		.out3_valid         (output_south_valid),              //      .valid
		.out3_ready         (output_south_ready),              //      .ready
		.out3_startofpacket (output_south_startofpacket),      //      .startofpacket
		.out3_endofpacket   (output_south_endofpacket),        //      .endofpacket
		.out3_empty         (output_south_empty),              //      .empty
		.out4_data          (output_east_data),                //  out4.data
		.out4_valid         (output_east_valid),               //      .valid
		.out4_ready         (output_east_ready),               //      .ready
		.out4_startofpacket (output_east_startofpacket),       //      .startofpacket
		.out4_endofpacket   (output_east_endofpacket),         //      .endofpacket
		.out4_empty         (output_east_empty)                //      .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
